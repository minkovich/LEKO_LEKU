Library IEEE;
	use IEEE.std_logic_1164.all;
entity x25_11x is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A76: buffer std_logic
);
end x25_11x;

architecture x25_11x_behav of x25_11x is
signal a1a,a2a,a3a,a4a,a5a,a6a,a7a,a8a,a9a,a10a,a11a,a12a,a13a,a14a,a15a,a16a,a17a,a18a,a19a,a20a,a21a,a22a,a23a,a24a,a25a,a26a,a27a,a28a,a29a,a30a,a31a,a32a,a33a,a34a,a35a,a36a,a37a,a38a,a39a,a40a,a41a,a42a,a43a,a44a,a45a,a46a,a47a,a48a,a49a,a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a159a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a172a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a251a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a313a,a314a,a315a,a316a,a317a,a318a,a319a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a353a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a405a,a406a,a407a,a408a,a409a,a410a,a411a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a456a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a537a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a551a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a655a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a735a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a807a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a838a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a,a854a,a855a,a856a,a857a,a858a,a859a,a860a,a861a,a862a,a863a,a864a,a865a,a866a,a867a,a868a,a869a,a870a,a871a,a872a,a873a,a874a,a875a,a876a,a877a,a878a,a879a,a880a,a881a,a882a,a883a,a884a,a885a,a886a,a887a,a888a,a889a,a890a,a891a,a892a,a893a,a894a,a895a,a896a,a897a,a898a,a899a,a900a,a901a,a902a,a903a,a904a,a905a,a906a,a907a,a908a,a909a,a910a,a911a,a912a,a913a,a914a,a915a,a916a,a917a,a918a,a919a,a920a,a921a,a922a,a923a,a924a,a925a,a926a,a927a,a928a,a929a,a930a,a931a,a932a,a933a,a934a,a935a,a936a,a937a,a938a,a939a,a940a,a941a,a942a,a943a,a944a,a945a,a946a,a947a,a948a,a949a,a950a,a951a,a952a,a953a,a954a,a955a,a956a,a957a,a958a,a959a,a960a,a961a,a962a,a963a,a964a,a965a,a966a,a967a,a968a,a969a,a970a,a971a,a972a,a973a,a974a,a975a,a976a,a977a,a978a,a979a,a980a,a981a,a982a,a983a,a984a,a985a,a986a,a987a,a988a,a989a,a990a,a991a,a992a,a993a,a994a,a995a,a996a,a997a,a998a,a999a,a1000a,a1001a,a1002a,a1003a,a1004a,a1005a,a1006a,a1007a,a1008a,a1009a,a1010a,a1011a,a1012a,a1013a,a1014a,a1015a,a1016a,a1017a,a1018a,a1019a,a1020a,a1021a,a1022a,a1023a,a1024a,a1025a,a1026a,a1027a,a1028a,a1029a,a1030a,a1031a,a1032a,a1033a,a1034a,a1035a,a1036a,a1037a,a1038a,a1039a,a1040a,a1041a,a1042a,a1043a,a1044a,a1045a,a1046a,a1047a,a1048a,a1049a,a1050a,a1051a,a1052a,a1053a,a1054a,a1055a,a1056a,a1057a,a1058a,a1059a,a1060a,a1061a,a1062a,a1063a,a1064a,a1065a,a1066a,a1067a,a1068a,a1069a,a1070a,a1071a,a1072a,a1073a,a1074a,a1075a,a1076a,a1077a,a1078a,a1079a,a1080a,a1081a,a1082a,a1083a,a1084a,a1085a,a1086a,a1087a,a1088a,a1089a,a1090a,a1091a,a1092a,a1093a,a1094a,a1095a,a1096a,a1097a,a1098a,a1099a,a1100a,a1101a,a1102a,a1103a,a1104a,a1105a,a1106a,a1107a,a1108a,a1109a,a1110a,a1111a,a1112a,a1113a,a1114a,a1115a,a1116a,a1117a,a1118a,a1119a,a1120a,a1121a,a1122a,a1123a,a1124a,a1125a,a1126a,a1127a,a1128a,a1129a,a1130a,a1131a,a1132a,a1133a,a1134a,a1135a,a1136a,a1137a,a1138a,a1139a,a1140a,a1141a,a1142a,a1143a,a1144a,a1145a,a1146a,a1147a,a1148a,a1149a,a1150a,a1151a,a1152a,a1153a,a1154a,a1155a,a1156a,a1157a,a1158a,a1159a,a1160a,a1161a,a1162a,a1163a,a1164a,a1165a,a1166a,a1167a,a1168a,a1169a,a1170a,a1171a,a1172a,a1173a,a1174a,a1175a,a1176a,a1177a,a1178a,a1179a,a1180a,a1181a,a1182a,a1183a,a1184a,a1185a,a1186a,a1187a,a1188a,a1189a,a1190a,a1191a,a1192a,a1193a,a1194a,a1195a,a1196a,a1197a,a1198a,a1199a,a1200a,a1201a,a1202a,a1203a,a1204a,a1205a,a1206a,a1207a,a1208a,a1209a,a1210a,a1211a,a1212a,a1213a,a1214a,a1215a,a1216a,a1217a,a1218a,a1219a,a1220a,a1221a,a1222a,a1223a,a1224a,a1225a,a1226a,a1227a,a1228a,a1229a,a1230a,a1231a,a1232a,a1233a,a1234a,a1235a,a1236a,a1237a,a1238a,a1239a,a1240a,a1241a,a1242a,a1243a,a1244a,a1245a,a1246a,a1247a,a1248a,a1249a,a1250a,a1251a,a1252a,a1253a,a1254a,a1255a,a1256a,a1257a,a1258a,a1259a,a1260a,a1261a,a1262a,a1263a,a1264a,a1265a,a1266a,a1267a,a1268a,a1269a,a1270a,a1271a,a1272a,a1273a,a1274a,a1275a,a1276a,a1277a,a1278a,a1279a,a1280a,a1281a,a1282a,a1283a,a1284a,a1285a,a1286a,a1287a,a1288a,a1289a,a1290a,a1291a,a1292a,a1293a,a1294a,a1295a,a1296a,a1297a,a1298a,a1299a,a1300a,a1301a,a1302a,a1303a,a1304a,a1305a,a1306a,a1307a,a1308a,a1309a,a1310a,a1311a,a1312a,a1313a,a1314a,a1315a,a1316a,a1317a,a1318a,a1319a,a1320a,a1321a,a1322a,a1323a,a1324a,a1325a,a1326a,a1327a,a1328a,a1329a,a1330a,a1331a,a1332a,a1333a,a1334a,a1335a,a1336a,a1337a,a1338a,a1339a,a1340a,a1341a,a1342a,a1343a,a1344a,a1345a,a1346a,a1347a,a1348a,a1349a,a1350a,a1351a,a1352a,a1353a,a1354a,a1355a,a1356a,a1357a,a1358a,a1359a,a1360a,a1361a,a1362a,a1363a,a1364a,a1365a,a1366a,a1367a,a1368a,a1369a,a1370a,a1371a,a1372a,a1373a,a1374a,a1375a,a1376a,a1377a,a1378a,a1379a,a1380a,a1381a,a1382a,a1383a,a1384a,a1385a,a1386a,a1387a,a1388a,a1389a,a1390a,a1391a,a1392a,a1393a,a1394a,a1395a,a1396a,a1397a,a1398a,a1399a,a1400a,a1401a,a1402a,a1403a,a1404a,a1405a,a1406a,a1407a,a1408a,a1409a,a1410a,a1411a,a1412a,a1413a,a1414a,a1415a,a1416a,a1417a,a1418a,a1419a,a1420a,a1421a,a1422a,a1423a,a1424a,a1425a,a1426a,a1427a,a1428a,a1429a,a1430a,a1431a,a1432a,a1433a,a1434a,a1435a,a1436a,a1437a,a1438a,a1439a,a1440a,a1441a,a1442a,a1443a,a1444a,a1445a,a1446a,a1447a,a1448a,a1449a,a1450a,a1451a,a1452a,a1453a,a1454a,a1455a,a1456a,a1457a,a1458a,a1459a,a1460a,a1461a,a1462a,a1463a,a1464a,a1465a,a1466a,a1467a,a1468a,a1469a,a1470a,a1471a,a1472a,a1473a,a1474a,a1475a,a1476a,a1477a,a1478a,a1479a,a1480a,a1481a,a1482a,a1483a,a1484a,a1485a,a1486a,a1487a,a1488a,a1489a,a1490a,a1491a,a1492a,a1493a,a1494a,a1495a,a1496a,a1497a,a1498a,a1499a,a1500a,a1501a,a1502a,a1503a,a1504a,a1505a,a1506a,a1507a,a1508a,a1509a,a1510a,a1511a,a1512a,a1513a,a1514a,a1515a,a1516a,a1517a,a1518a,a1519a,a1520a,a1521a,a1522a,a1523a,a1524a,a1525a,a1526a,a1527a,a1528a,a1529a,a1530a,a1531a,a1532a,a1533a,a1534a,a1535a,a1536a,a1537a,a1538a,a1539a,a1540a,a1541a,a1542a,a1543a,a1544a,a1545a,a1546a,a1547a,a1548a,a1549a,a1550a,a1551a,a1552a,a1553a,a1554a,a1555a,a1556a,a1557a,a1558a,a1559a,a1560a,a1561a,a1562a,a1563a,a1564a,a1565a,a1566a,a1567a,a1568a,a1569a,a1570a,a1571a,a1572a,a1573a,a1574a,a1575a,a1576a,a1577a,a1578a,a1579a,a1580a,a1581a,a1582a,a1583a,a1584a,a1585a,a1586a,a1587a,a1588a,a1589a,a1590a,a1591a,a1592a,a1593a,a1594a,a1595a,a1596a,a1597a,a1598a,a1599a,a1600a,a1601a,a1602a,a1603a,a1604a,a1605a,a1606a,a1607a,a1608a,a1609a,a1610a,a1611a,a1612a,a1613a,a1614a,a1615a,a1616a,a1617a,a1618a,a1619a,a1620a,a1621a,a1622a,a1623a,a1624a,a1625a,a1626a,a1627a,a1628a,a1629a,a1630a,a1631a,a1632a,a1633a,a1634a,a1635a,a1636a,a1637a,a1638a,a1639a,a1640a,a1641a,a1642a,a1643a,a1644a,a1645a,a1646a,a1647a,a1648a,a1649a,a1650a,a1651a,a1652a,a1653a,a1654a,a1655a,a1656a,a1657a,a1658a,a1659a,a1660a,a1661a,a1662a,a1663a,a1664a,a1665a,a1666a,a1667a,a1668a,a1669a,a1670a,a1671a,a1672a,a1673a,a1674a,a1675a,a1676a,a1677a,a1678a,a1679a,a1680a,a1681a,a1682a,a1683a,a1684a,a1685a,a1686a,a1687a,a1688a,a1689a,a1690a,a1691a,a1692a,a1693a,a1694a,a1695a,a1696a,a1697a,a1698a,a1699a,a1700a,a1701a,a1702a,a1703a,a1704a,a1705a,a1706a,a1707a,a1708a,a1709a,a1710a,a1711a,a1712a,a1713a,a1714a,a1715a,a1716a,a1717a,a1718a,a1719a,a1720a,a1721a,a1722a,a1723a,a1724a,a1725a,a1726a,a1727a,a1728a,a1729a,a1730a,a1731a,a1732a,a1733a,a1734a,a1735a,a1736a,a1737a,a1738a,a1739a,a1740a,a1741a,a1742a,a1743a,a1744a,a1745a,a1746a,a1747a,a1748a,a1749a,a1750a,a1751a,a1752a,a1753a,a1754a,a1755a,a1756a,a1757a,a1758a,a1759a,a1760a,a1761a,a1762a,a1763a,a1764a,a1765a,a1766a,a1767a,a1768a,a1769a,a1770a,a1771a,a1772a,a1773a,a1774a,a1775a,a1776a,a1777a,a1778a,a1779a,a1780a,a1781a,a1782a,a1783a,a1784a,a1785a,a1786a,a1787a,a1788a,a1789a,a1790a,a1791a,a1792a,a1793a,a1794a,a1795a,a1796a,a1797a,a1798a,a1799a,a1800a,a1801a,a1802a,a1803a,a1804a,a1805a,a1806a,a1807a,a1808a,a1809a,a1810a,a1811a,a1812a,a1813a,a1814a,a1815a,a1816a,a1817a,a1818a,a1819a,a1820a,a1821a,a1822a,a1823a,a1824a,a1825a,a1826a,a1827a,a1828a,a1829a,a1830a,a1831a,a1832a,a1833a,a1834a,a1835a,a1836a,a1837a,a1838a,a1839a,a1840a,a1841a,a1842a,a1843a,a1844a,a1845a,a1846a,a1847a,a1848a,a1849a,a1850a,a1851a,a1852a,a1853a,a1854a,a1855a,a1856a,a1857a,a1858a,a1859a,a1860a,a1861a,a1862a,a1863a,a1864a,a1865a,a1866a,a1867a,a1868a,a1869a,a1870a,a1871a,a1872a,a1873a,a1874a,a1875a,a1876a,a1877a,a1878a,a1879a,a1880a,a1881a,a1882a,a1883a,a1884a,a1885a,a1886a,a1887a,a1888a,a1889a,a1890a,a1891a,a1892a,a1893a,a1894a,a1895a,a1896a,a1897a,a1898a,a1899a,a1900a,a1901a,a1902a,a1903a,a1904a,a1905a,a1906a,a1907a,a1908a,a1909a,a1910a,a1911a,a1912a,a1913a,a1914a,a1915a,a1916a,a1917a,a1918a,a1919a,a1920a,a1921a,a1922a,a1923a,a1924a,a1925a,a1926a,a1927a,a1928a,a1929a,a1930a,a1931a,a1932a,a1933a,a1934a,a1935a,a1936a,a1937a,a1938a,a1939a,a1940a,a1941a,a1942a,a1943a,a1944a,a1945a,a1946a,a1947a,a1948a,a1949a,a1950a,a1951a,a1952a,a1953a,a1954a,a1955a,a1956a,a1957a,a1958a,a1959a,a1960a,a1961a,a1962a,a1963a,a1964a,a1965a,a1966a,a1967a,a1968a,a1969a,a1970a,a1971a,a1972a,a1973a,a1974a,a1975a,a1976a,a1977a,a1978a,a1979a,a1980a,a1981a,a1982a,a1983a,a1984a,a1985a,a1986a,a1987a,a1988a,a1989a,a1990a,a1991a,a1992a,a1993a,a1994a,a1995a,a1996a,a1997a,a1998a,a1999a,a2000a,a2001a,a2002a,a2003a,a2004a,a2005a,a2006a,a2007a,a2008a,a2009a,a2010a,a2011a,a2012a,a2013a,a2014a,a2015a,a2016a,a2017a,a2018a,a2019a,a2020a,a2021a,a2022a,a2023a,a2024a,a2025a,a2026a,a2027a,a2028a,a2029a,a2030a,a2031a,a2032a,a2033a,a2034a,a2035a,a2036a,a2037a,a2038a,a2039a,a2040a,a2041a,a2042a,a2043a,a2044a,a2045a,a2046a,a2047a,a2048a,a2049a,a2050a,a2051a,a2052a,a2053a,a2054a,a2055a,a2056a,a2057a,a2058a,a2059a,a2060a,a2061a,a2062a,a2063a,a2064a,a2065a,a2066a,a2067a,a2068a,a2069a,a2070a,a2071a,a2072a,a2073a,a2074a,a2075a,a2076a,a2077a,a2078a,a2079a,a2080a,a2081a,a2082a,a2083a,a2084a,a2085a,a2086a,a2087a,a2088a,a2089a,a2090a,a2091a,a2092a,a2093a,a2094a,a2095a,a2096a,a2097a,a2098a,a2099a,a2100a,a2101a,a2102a,a2103a,a2104a,a2105a,a2106a,a2107a,a2108a,a2109a,a2110a,a2111a,a2112a,a2113a,a2114a,a2115a,a2116a,a2117a,a2118a,a2119a,a2120a,a2121a,a2122a,a2123a,a2124a,a2125a,a2126a,a2127a,a2128a,a2129a,a2130a,a2131a,a2132a,a2133a,a2134a,a2135a,a2136a,a2137a,a2138a,a2139a,a2140a,a2141a,a2142a,a2143a,a2144a,a2145a,a2146a,a2147a,a2148a,a2149a,a2150a,a2151a,a2152a,a2153a,a2154a,a2155a,a2156a,a2157a,a2158a,a2159a,a2160a,a2161a,a2162a,a2163a,a2164a,a2165a,a2166a,a2167a,a2168a,a2169a,a2170a,a2171a,a2172a,a2173a,a2174a,a2175a,a2176a,a2177a,a2178a,a2179a,a2180a,a2181a,a2182a,a2183a,a2184a,a2185a,a2186a,a2187a,a2188a,a2189a,a2190a,a2191a,a2192a,a2193a,a2194a,a2195a,a2196a,a2197a,a2198a,a2199a,a2200a,a2201a,a2202a,a2203a,a2204a,a2205a,a2206a,a2207a,a2208a,a2209a,a2210a,a2211a,a2212a,a2213a,a2214a,a2215a,a2216a,a2217a,a2218a,a2219a,a2220a,a2221a,a2222a,a2223a,a2224a,a2225a,a2226a,a2227a,a2228a,a2229a,a2230a,a2231a,a2232a,a2233a,a2234a,a2235a,a2236a,a2237a,a2238a,a2239a,a2240a,a2241a,a2242a,a2243a,a2244a,a2245a,a2246a,a2247a,a2248a,a2249a,a2250a,a2251a,a2252a,a2253a,a2254a,a2255a,a2256a,a2257a,a2258a,a2259a,a2260a,a2261a,a2262a,a2263a,a2264a,a2265a,a2266a,a2267a,a2268a,a2269a,a2270a,a2271a,a2272a,a2273a,a2274a,a2275a,a2276a,a2277a,a2278a,a2279a,a2280a,a2281a,a2282a,a2283a,a2284a,a2285a,a2286a,a2287a,a2288a,a2289a,a2290a,a2291a,a2292a,a2293a,a2294a,a2295a,a2296a,a2297a,a2298a,a2299a,a2300a,a2301a,a2302a,a2303a,a2304a,a2305a,a2306a,a2307a,a2308a,a2309a,a2310a,a2313a,a2316a,a2317a,a2320a,a2324a,a2325a,a2326a,a2327a,a2330a,a2333a,a2334a,a2337a,a2341a,a2342a,a2343a,a2344a,a2345a,a2348a,a2351a,a2352a,a2355a,a2359a,a2360a,a2361a,a2362a,a2365a,a2368a,a2369a,a2372a,a2376a,a2377a,a2378a,a2379a,a2380a,a2381a,a2384a,a2387a,a2388a,a2391a,a2395a,a2396a,a2397a,a2398a,a2401a,a2404a,a2405a,a2408a,a2412a,a2413a,a2414a,a2415a,a2416a,a2419a,a2422a,a2423a,a2426a,a2430a,a2431a,a2432a,a2433a,a2436a,a2439a,a2440a,a2443a,a2447a,a2448a,a2449a,a2450a,a2451a,a2452a,a2453a,a2456a,a2459a,a2460a,a2463a,a2467a,a2468a,a2469a,a2470a,a2473a,a2476a,a2477a,a2480a,a2484a,a2485a,a2486a,a2487a,a2488a,a2491a,a2494a,a2495a,a2498a,a2502a,a2503a,a2504a,a2505a,a2508a,a2511a,a2512a,a2515a,a2519a,a2520a,a2521a,a2522a,a2523a,a2524a,a2527a,a2530a,a2531a,a2534a,a2538a,a2539a,a2540a,a2541a,a2544a,a2547a,a2548a,a2551a,a2555a,a2556a,a2557a,a2558a,a2559a,a2562a,a2565a,a2566a,a2569a,a2573a,a2574a,a2575a,a2576a,a2579a,a2582a,a2583a,a2586a,a2590a,a2591a,a2592a,a2593a,a2594a,a2595a,a2596a,a2597a,a2600a,a2603a,a2604a,a2607a,a2611a,a2612a,a2613a,a2614a,a2617a,a2620a,a2621a,a2624a,a2628a,a2629a,a2630a,a2631a,a2632a,a2635a,a2638a,a2639a,a2642a,a2646a,a2647a,a2648a,a2649a,a2652a,a2655a,a2656a,a2659a,a2663a,a2664a,a2665a,a2666a,a2667a,a2668a,a2671a,a2674a,a2675a,a2678a,a2682a,a2683a,a2684a,a2685a,a2688a,a2691a,a2692a,a2695a,a2699a,a2700a,a2701a,a2702a,a2703a,a2706a,a2709a,a2710a,a2713a,a2717a,a2718a,a2719a,a2720a,a2723a,a2726a,a2727a,a2730a,a2734a,a2735a,a2736a,a2737a,a2738a,a2739a,a2740a,a2743a,a2746a,a2747a,a2750a,a2754a,a2755a,a2756a,a2757a,a2760a,a2763a,a2764a,a2767a,a2771a,a2772a,a2773a,a2774a,a2775a,a2778a,a2781a,a2782a,a2785a,a2789a,a2790a,a2791a,a2792a,a2795a,a2798a,a2799a,a2802a,a2806a,a2807a,a2808a,a2809a,a2810a,a2811a,a2814a,a2817a,a2818a,a2821a,a2825a,a2826a,a2827a,a2828a,a2831a,a2834a,a2835a,a2838a,a2842a,a2843a,a2844a,a2845a,a2846a,a2849a,a2852a,a2853a,a2856a,a2860a,a2861a,a2862a,a2863a,a2866a,a2869a,a2870a,a2873a,a2877a,a2878a,a2879a,a2880a,a2881a,a2882a,a2883a,a2884a,a2885a,a2888a,a2891a,a2892a,a2895a,a2899a,a2900a,a2901a,a2902a,a2905a,a2908a,a2909a,a2912a,a2916a,a2917a,a2918a,a2919a,a2920a,a2923a,a2926a,a2927a,a2930a,a2934a,a2935a,a2936a,a2937a,a2940a,a2943a,a2944a,a2947a,a2951a,a2952a,a2953a,a2954a,a2955a,a2956a,a2959a,a2962a,a2963a,a2966a,a2970a,a2971a,a2972a,a2973a,a2976a,a2979a,a2980a,a2983a,a2987a,a2988a,a2989a,a2990a,a2991a,a2994a,a2997a,a2998a,a3001a,a3005a,a3006a,a3007a,a3008a,a3011a,a3014a,a3015a,a3018a,a3022a,a3023a,a3024a,a3025a,a3026a,a3027a,a3028a,a3031a,a3034a,a3035a,a3038a,a3042a,a3043a,a3044a,a3045a,a3048a,a3051a,a3052a,a3055a,a3059a,a3060a,a3061a,a3062a,a3063a,a3066a,a3069a,a3070a,a3073a,a3077a,a3078a,a3079a,a3080a,a3083a,a3086a,a3087a,a3090a,a3094a,a3095a,a3096a,a3097a,a3098a,a3099a,a3102a,a3105a,a3106a,a3109a,a3113a,a3114a,a3115a,a3116a,a3119a,a3122a,a3123a,a3126a,a3130a,a3131a,a3132a,a3133a,a3134a,a3137a,a3140a,a3141a,a3144a,a3148a,a3149a,a3150a,a3151a,a3154a,a3157a,a3158a,a3161a,a3165a,a3166a,a3167a,a3168a,a3169a,a3170a,a3171a,a3172a,a3175a,a3178a,a3179a,a3182a,a3186a,a3187a,a3188a,a3189a,a3192a,a3195a,a3196a,a3199a,a3203a,a3204a,a3205a,a3206a,a3207a,a3210a,a3213a,a3214a,a3217a,a3221a,a3222a,a3223a,a3224a,a3227a,a3230a,a3231a,a3234a,a3238a,a3239a,a3240a,a3241a,a3242a,a3243a,a3246a,a3249a,a3250a,a3253a,a3257a,a3258a,a3259a,a3260a,a3263a,a3266a,a3267a,a3270a,a3274a,a3275a,a3276a,a3277a,a3278a,a3281a,a3284a,a3285a,a3288a,a3292a,a3293a,a3294a,a3295a,a3298a,a3301a,a3302a,a3305a,a3309a,a3310a,a3311a,a3312a,a3313a,a3314a,a3315a,a3318a,a3321a,a3322a,a3325a,a3329a,a3330a,a3331a,a3332a,a3335a,a3338a,a3339a,a3342a,a3346a,a3347a,a3348a,a3349a,a3350a,a3353a,a3356a,a3357a,a3360a,a3364a,a3365a,a3366a,a3367a,a3370a,a3373a,a3374a,a3377a,a3381a,a3382a,a3383a,a3384a,a3385a,a3386a,a3389a,a3392a,a3393a,a3396a,a3400a,a3401a,a3402a,a3403a,a3406a,a3409a,a3410a,a3413a,a3417a,a3418a,a3419a,a3420a,a3421a,a3424a,a3427a,a3428a,a3431a,a3435a,a3436a,a3437a,a3438a,a3441a,a3445a,a3446a,a3447a,a3450a,a3454a,a3455a,a3456a,a3457a,a3458a,a3459a,a3460a,a3461a,a3462a,a3463a,a3466a,a3469a,a3470a,a3473a,a3477a,a3478a,a3479a,a3480a,a3483a,a3486a,a3487a,a3490a,a3494a,a3495a,a3496a,a3497a,a3498a,a3501a,a3504a,a3505a,a3508a,a3512a,a3513a,a3514a,a3515a,a3518a,a3521a,a3522a,a3525a,a3529a,a3530a,a3531a,a3532a,a3533a,a3534a,a3537a,a3540a,a3541a,a3544a,a3548a,a3549a,a3550a,a3551a,a3554a,a3557a,a3558a,a3561a,a3565a,a3566a,a3567a,a3568a,a3569a,a3572a,a3575a,a3576a,a3579a,a3583a,a3584a,a3585a,a3586a,a3589a,a3592a,a3593a,a3596a,a3600a,a3601a,a3602a,a3603a,a3604a,a3605a,a3606a,a3609a,a3612a,a3613a,a3616a,a3620a,a3621a,a3622a,a3623a,a3626a,a3629a,a3630a,a3633a,a3637a,a3638a,a3639a,a3640a,a3641a,a3644a,a3647a,a3648a,a3651a,a3655a,a3656a,a3657a,a3658a,a3661a,a3664a,a3665a,a3668a,a3672a,a3673a,a3674a,a3675a,a3676a,a3677a,a3680a,a3683a,a3684a,a3687a,a3691a,a3692a,a3693a,a3694a,a3697a,a3700a,a3701a,a3704a,a3708a,a3709a,a3710a,a3711a,a3712a,a3715a,a3718a,a3719a,a3722a,a3726a,a3727a,a3728a,a3729a,a3732a,a3735a,a3736a,a3739a,a3743a,a3744a,a3745a,a3746a,a3747a,a3748a,a3749a,a3750a,a3753a,a3756a,a3757a,a3760a,a3764a,a3765a,a3766a,a3767a,a3770a,a3773a,a3774a,a3777a,a3781a,a3782a,a3783a,a3784a,a3785a,a3788a,a3791a,a3792a,a3795a,a3799a,a3800a,a3801a,a3802a,a3805a,a3808a,a3809a,a3812a,a3816a,a3817a,a3818a,a3819a,a3820a,a3821a,a3824a,a3827a,a3828a,a3831a,a3835a,a3836a,a3837a,a3838a,a3841a,a3844a,a3845a,a3848a,a3852a,a3853a,a3854a,a3855a,a3856a,a3859a,a3862a,a3863a,a3866a,a3870a,a3871a,a3872a,a3873a,a3876a,a3879a,a3880a,a3883a,a3887a,a3888a,a3889a,a3890a,a3891a,a3892a,a3893a,a3896a,a3899a,a3900a,a3903a,a3907a,a3908a,a3909a,a3910a,a3913a,a3916a,a3917a,a3920a,a3924a,a3925a,a3926a,a3927a,a3928a,a3931a,a3934a,a3935a,a3938a,a3942a,a3943a,a3944a,a3945a,a3948a,a3951a,a3952a,a3955a,a3959a,a3960a,a3961a,a3962a,a3963a,a3964a,a3967a,a3970a,a3971a,a3974a,a3978a,a3979a,a3980a,a3981a,a3984a,a3987a,a3988a,a3991a,a3995a,a3996a,a3997a,a3998a,a3999a,a4002a,a4005a,a4006a,a4009a,a4013a,a4014a,a4015a,a4016a,a4019a,a4023a,a4024a,a4025a,a4028a,a4032a,a4033a,a4034a,a4035a,a4036a,a4037a,a4038a,a4039a,a4040a,a4043a,a4046a,a4047a,a4050a,a4054a,a4055a,a4056a,a4057a,a4060a,a4063a,a4064a,a4067a,a4071a,a4072a,a4073a,a4074a,a4075a,a4078a,a4081a,a4082a,a4085a,a4089a,a4090a,a4091a,a4092a,a4095a,a4098a,a4099a,a4102a,a4106a,a4107a,a4108a,a4109a,a4110a,a4111a,a4114a,a4117a,a4118a,a4121a,a4125a,a4126a,a4127a,a4128a,a4131a,a4134a,a4135a,a4138a,a4142a,a4143a,a4144a,a4145a,a4146a,a4149a,a4152a,a4153a,a4156a,a4160a,a4161a,a4162a,a4163a,a4166a,a4169a,a4170a,a4173a,a4177a,a4178a,a4179a,a4180a,a4181a,a4182a,a4183a,a4186a,a4189a,a4190a,a4193a,a4197a,a4198a,a4199a,a4200a,a4203a,a4206a,a4207a,a4210a,a4214a,a4215a,a4216a,a4217a,a4218a,a4221a,a4224a,a4225a,a4228a,a4232a,a4233a,a4234a,a4235a,a4238a,a4241a,a4242a,a4245a,a4249a,a4250a,a4251a,a4252a,a4253a,a4254a,a4257a,a4260a,a4261a,a4264a,a4268a,a4269a,a4270a,a4271a,a4274a,a4277a,a4278a,a4281a,a4285a,a4286a,a4287a,a4288a,a4289a,a4292a,a4295a,a4296a,a4299a,a4303a,a4304a,a4305a,a4306a,a4309a,a4312a,a4313a,a4316a,a4320a,a4321a,a4322a,a4323a,a4324a,a4325a,a4326a,a4327a,a4330a,a4333a,a4334a,a4337a,a4341a,a4342a,a4343a,a4344a,a4347a,a4350a,a4351a,a4354a,a4358a,a4359a,a4360a,a4361a,a4362a,a4365a,a4368a,a4369a,a4372a,a4376a,a4377a,a4378a,a4379a,a4382a,a4385a,a4386a,a4389a,a4393a,a4394a,a4395a,a4396a,a4397a,a4398a,a4401a,a4404a,a4405a,a4408a,a4412a,a4413a,a4414a,a4415a,a4418a,a4421a,a4422a,a4425a,a4429a,a4430a,a4431a,a4432a,a4433a,a4436a,a4439a,a4440a,a4443a,a4447a,a4448a,a4449a,a4450a,a4453a,a4456a,a4457a,a4460a,a4464a,a4465a,a4466a,a4467a,a4468a,a4469a,a4470a,a4473a,a4476a,a4477a,a4480a,a4484a,a4485a,a4486a,a4487a,a4490a,a4493a,a4494a,a4497a,a4501a,a4502a,a4503a,a4504a,a4505a,a4508a,a4511a,a4512a,a4515a,a4519a,a4520a,a4521a,a4522a,a4525a,a4528a,a4529a,a4532a,a4536a,a4537a,a4538a,a4539a,a4540a,a4541a,a4544a,a4547a,a4548a,a4551a,a4555a,a4556a,a4557a,a4558a,a4561a,a4564a,a4565a,a4568a,a4572a,a4573a,a4574a,a4575a,a4576a,a4579a,a4582a,a4583a,a4586a,a4590a,a4591a,a4592a,a4593a,a4596a,a4600a,a4601a,a4602a,a4605a,a4609a,a4610a,a4611a,a4612a,a4613a,a4614a,a4615a,a4616a,a4617a,a4618a,a4619a,a4622a,a4625a,a4626a,a4629a,a4633a,a4634a,a4635a,a4636a,a4639a,a4642a,a4643a,a4646a,a4650a,a4651a,a4652a,a4653a,a4654a,a4657a,a4660a,a4661a,a4664a,a4668a,a4669a,a4670a,a4671a,a4674a,a4677a,a4678a,a4681a,a4685a,a4686a,a4687a,a4688a,a4689a,a4690a,a4693a,a4696a,a4697a,a4700a,a4704a,a4705a,a4706a,a4707a,a4710a,a4713a,a4714a,a4717a,a4721a,a4722a,a4723a,a4724a,a4725a,a4728a,a4731a,a4732a,a4735a,a4739a,a4740a,a4741a,a4742a,a4745a,a4748a,a4749a,a4752a,a4756a,a4757a,a4758a,a4759a,a4760a,a4761a,a4762a,a4765a,a4768a,a4769a,a4772a,a4776a,a4777a,a4778a,a4779a,a4782a,a4785a,a4786a,a4789a,a4793a,a4794a,a4795a,a4796a,a4797a,a4800a,a4803a,a4804a,a4807a,a4811a,a4812a,a4813a,a4814a,a4817a,a4820a,a4821a,a4824a,a4828a,a4829a,a4830a,a4831a,a4832a,a4833a,a4836a,a4839a,a4840a,a4843a,a4847a,a4848a,a4849a,a4850a,a4853a,a4856a,a4857a,a4860a,a4864a,a4865a,a4866a,a4867a,a4868a,a4871a,a4874a,a4875a,a4878a,a4882a,a4883a,a4884a,a4885a,a4888a,a4891a,a4892a,a4895a,a4899a,a4900a,a4901a,a4902a,a4903a,a4904a,a4905a,a4906a,a4909a,a4912a,a4913a,a4916a,a4920a,a4921a,a4922a,a4923a,a4926a,a4929a,a4930a,a4933a,a4937a,a4938a,a4939a,a4940a,a4941a,a4944a,a4947a,a4948a,a4951a,a4955a,a4956a,a4957a,a4958a,a4961a,a4964a,a4965a,a4968a,a4972a,a4973a,a4974a,a4975a,a4976a,a4977a,a4980a,a4983a,a4984a,a4987a,a4991a,a4992a,a4993a,a4994a,a4997a,a5000a,a5001a,a5004a,a5008a,a5009a,a5010a,a5011a,a5012a,a5015a,a5018a,a5019a,a5022a,a5026a,a5027a,a5028a,a5029a,a5032a,a5035a,a5036a,a5039a,a5043a,a5044a,a5045a,a5046a,a5047a,a5048a,a5049a,a5052a,a5055a,a5056a,a5059a,a5063a,a5064a,a5065a,a5066a,a5069a,a5072a,a5073a,a5076a,a5080a,a5081a,a5082a,a5083a,a5084a,a5087a,a5090a,a5091a,a5094a,a5098a,a5099a,a5100a,a5101a,a5104a,a5107a,a5108a,a5111a,a5115a,a5116a,a5117a,a5118a,a5119a,a5120a,a5123a,a5126a,a5127a,a5130a,a5134a,a5135a,a5136a,a5137a,a5140a,a5143a,a5144a,a5147a,a5151a,a5152a,a5153a,a5154a,a5155a,a5158a,a5161a,a5162a,a5165a,a5169a,a5170a,a5171a,a5172a,a5175a,a5178a,a5179a,a5182a,a5186a,a5187a,a5188a,a5189a,a5190a,a5191a,a5192a,a5193a,a5194a,a5197a,a5200a,a5201a,a5204a,a5208a,a5209a,a5210a,a5211a,a5214a,a5217a,a5218a,a5221a,a5225a,a5226a,a5227a,a5228a,a5229a,a5232a,a5235a,a5236a,a5239a,a5243a,a5244a,a5245a,a5246a,a5249a,a5252a,a5253a,a5256a,a5260a,a5261a,a5262a,a5263a,a5264a,a5265a,a5268a,a5271a,a5272a,a5275a,a5279a,a5280a,a5281a,a5282a,a5285a,a5288a,a5289a,a5292a,a5296a,a5297a,a5298a,a5299a,a5300a,a5303a,a5306a,a5307a,a5310a,a5314a,a5315a,a5316a,a5317a,a5320a,a5323a,a5324a,a5327a,a5331a,a5332a,a5333a,a5334a,a5335a,a5336a,a5337a,a5340a,a5343a,a5344a,a5347a,a5351a,a5352a,a5353a,a5354a,a5357a,a5360a,a5361a,a5364a,a5368a,a5369a,a5370a,a5371a,a5372a,a5375a,a5378a,a5379a,a5382a,a5386a,a5387a,a5388a,a5389a,a5392a,a5395a,a5396a,a5399a,a5403a,a5404a,a5405a,a5406a,a5407a,a5408a,a5411a,a5414a,a5415a,a5418a,a5422a,a5423a,a5424a,a5425a,a5428a,a5431a,a5432a,a5435a,a5439a,a5440a,a5441a,a5442a,a5443a,a5446a,a5449a,a5450a,a5453a,a5457a,a5458a,a5459a,a5460a,a5463a,a5466a,a5467a,a5470a,a5474a,a5475a,a5476a,a5477a,a5478a,a5479a,a5480a,a5481a,a5484a,a5487a,a5488a,a5491a,a5495a,a5496a,a5497a,a5498a,a5501a,a5504a,a5505a,a5508a,a5512a,a5513a,a5514a,a5515a,a5516a,a5519a,a5522a,a5523a,a5526a,a5530a,a5531a,a5532a,a5533a,a5536a,a5539a,a5540a,a5543a,a5547a,a5548a,a5549a,a5550a,a5551a,a5552a,a5555a,a5558a,a5559a,a5562a,a5566a,a5567a,a5568a,a5569a,a5572a,a5575a,a5576a,a5579a,a5583a,a5584a,a5585a,a5586a,a5587a,a5590a,a5593a,a5594a,a5597a,a5601a,a5602a,a5603a,a5604a,a5607a,a5610a,a5611a,a5614a,a5618a,a5619a,a5620a,a5621a,a5622a,a5623a,a5624a,a5627a,a5630a,a5631a,a5634a,a5638a,a5639a,a5640a,a5641a,a5644a,a5647a,a5648a,a5651a,a5655a,a5656a,a5657a,a5658a,a5659a,a5662a,a5665a,a5666a,a5669a,a5673a,a5674a,a5675a,a5676a,a5679a,a5682a,a5683a,a5686a,a5690a,a5691a,a5692a,a5693a,a5694a,a5695a,a5698a,a5701a,a5702a,a5705a,a5709a,a5710a,a5711a,a5712a,a5715a,a5718a,a5719a,a5722a,a5726a,a5727a,a5728a,a5729a,a5730a,a5733a,a5736a,a5737a,a5740a,a5744a,a5745a,a5746a,a5747a,a5750a,a5754a,a5755a,a5756a,a5759a,a5763a,a5764a,a5765a,a5766a,a5767a,a5768a,a5769a,a5770a,a5771a,a5772a,a5775a,a5778a,a5779a,a5782a,a5786a,a5787a,a5788a,a5789a,a5792a,a5795a,a5796a,a5799a,a5803a,a5804a,a5805a,a5806a,a5807a,a5810a,a5813a,a5814a,a5817a,a5821a,a5822a,a5823a,a5824a,a5827a,a5830a,a5831a,a5834a,a5838a,a5839a,a5840a,a5841a,a5842a,a5843a,a5846a,a5849a,a5850a,a5853a,a5857a,a5858a,a5859a,a5860a,a5863a,a5866a,a5867a,a5870a,a5874a,a5875a,a5876a,a5877a,a5878a,a5881a,a5884a,a5885a,a5888a,a5892a,a5893a,a5894a,a5895a,a5898a,a5901a,a5902a,a5905a,a5909a,a5910a,a5911a,a5912a,a5913a,a5914a,a5915a,a5918a,a5921a,a5922a,a5925a,a5929a,a5930a,a5931a,a5932a,a5935a,a5938a,a5939a,a5942a,a5946a,a5947a,a5948a,a5949a,a5950a,a5953a,a5956a,a5957a,a5960a,a5964a,a5965a,a5966a,a5967a,a5970a,a5973a,a5974a,a5977a,a5981a,a5982a,a5983a,a5984a,a5985a,a5986a,a5989a,a5992a,a5993a,a5996a,a6000a,a6001a,a6002a,a6003a,a6006a,a6009a,a6010a,a6013a,a6017a,a6018a,a6019a,a6020a,a6021a,a6024a,a6027a,a6028a,a6031a,a6035a,a6036a,a6037a,a6038a,a6041a,a6044a,a6045a,a6048a,a6052a,a6053a,a6054a,a6055a,a6056a,a6057a,a6058a,a6059a,a6062a,a6065a,a6066a,a6069a,a6073a,a6074a,a6075a,a6076a,a6079a,a6082a,a6083a,a6086a,a6090a,a6091a,a6092a,a6093a,a6094a,a6097a,a6100a,a6101a,a6104a,a6108a,a6109a,a6110a,a6111a,a6114a,a6117a,a6118a,a6121a,a6125a,a6126a,a6127a,a6128a,a6129a,a6130a,a6133a,a6136a,a6137a,a6140a,a6144a,a6145a,a6146a,a6147a,a6150a,a6153a,a6154a,a6157a,a6161a,a6162a,a6163a,a6164a,a6165a,a6168a,a6171a,a6172a,a6175a,a6179a,a6180a,a6181a,a6182a,a6185a,a6188a,a6189a,a6192a,a6196a,a6197a,a6198a,a6199a,a6200a,a6201a,a6202a,a6205a,a6208a,a6209a,a6212a,a6216a,a6217a,a6218a,a6219a,a6222a,a6225a,a6226a,a6229a,a6233a,a6234a,a6235a,a6236a,a6237a,a6240a,a6243a,a6244a,a6247a,a6251a,a6252a,a6253a,a6254a,a6257a,a6260a,a6261a,a6264a,a6268a,a6269a,a6270a,a6271a,a6272a,a6273a,a6276a,a6279a,a6280a,a6283a,a6287a,a6288a,a6289a,a6290a,a6293a,a6296a,a6297a,a6300a,a6304a,a6305a,a6306a,a6307a,a6308a,a6311a,a6314a,a6315a,a6318a,a6322a,a6323a,a6324a,a6325a,a6328a,a6332a,a6333a,a6334a,a6337a,a6341a,a6342a,a6343a,a6344a,a6345a,a6346a,a6347a,a6348a,a6349a,a6352a,a6355a,a6356a,a6359a,a6363a,a6364a,a6365a,a6366a,a6369a,a6372a,a6373a,a6376a,a6380a,a6381a,a6382a,a6383a,a6384a,a6387a,a6390a,a6391a,a6394a,a6398a,a6399a,a6400a,a6401a,a6404a,a6407a,a6408a,a6411a,a6415a,a6416a,a6417a,a6418a,a6419a,a6420a,a6423a,a6426a,a6427a,a6430a,a6434a,a6435a,a6436a,a6437a,a6440a,a6443a,a6444a,a6447a,a6451a,a6452a,a6453a,a6454a,a6455a,a6458a,a6461a,a6462a,a6465a,a6469a,a6470a,a6471a,a6472a,a6475a,a6478a,a6479a,a6482a,a6486a,a6487a,a6488a,a6489a,a6490a,a6491a,a6492a,a6495a,a6498a,a6499a,a6502a,a6506a,a6507a,a6508a,a6509a,a6512a,a6515a,a6516a,a6519a,a6523a,a6524a,a6525a,a6526a,a6527a,a6530a,a6533a,a6534a,a6537a,a6541a,a6542a,a6543a,a6544a,a6547a,a6550a,a6551a,a6554a,a6558a,a6559a,a6560a,a6561a,a6562a,a6563a,a6566a,a6569a,a6570a,a6573a,a6577a,a6578a,a6579a,a6580a,a6583a,a6586a,a6587a,a6590a,a6594a,a6595a,a6596a,a6597a,a6598a,a6601a,a6604a,a6605a,a6608a,a6612a,a6613a,a6614a,a6615a,a6618a,a6621a,a6622a,a6625a,a6629a,a6630a,a6631a,a6632a,a6633a,a6634a,a6635a,a6636a,a6639a,a6642a,a6643a,a6646a,a6650a,a6651a,a6652a,a6653a,a6656a,a6659a,a6660a,a6663a,a6667a,a6668a,a6669a,a6670a,a6671a,a6674a,a6677a,a6678a,a6681a,a6685a,a6686a,a6687a,a6688a,a6691a,a6694a,a6695a,a6698a,a6702a,a6703a,a6704a,a6705a,a6706a,a6707a,a6710a,a6713a,a6714a,a6717a,a6721a,a6722a,a6723a,a6724a,a6727a,a6730a,a6731a,a6734a,a6738a,a6739a,a6740a,a6741a,a6742a,a6745a,a6748a,a6749a,a6752a,a6756a,a6757a,a6758a,a6759a,a6762a,a6765a,a6766a,a6769a,a6773a,a6774a,a6775a,a6776a,a6777a,a6778a,a6779a,a6782a,a6785a,a6786a,a6789a,a6793a,a6794a,a6795a,a6796a,a6799a,a6802a,a6803a,a6806a,a6810a,a6811a,a6812a,a6813a,a6814a,a6817a,a6820a,a6821a,a6824a,a6828a,a6829a,a6830a,a6831a,a6834a,a6837a,a6838a,a6841a,a6845a,a6846a,a6847a,a6848a,a6849a,a6850a,a6853a,a6856a,a6857a,a6860a,a6864a,a6865a,a6866a,a6867a,a6870a,a6873a,a6874a,a6877a,a6881a,a6882a,a6883a,a6884a,a6885a,a6888a,a6891a,a6892a,a6895a,a6899a,a6900a,a6901a,a6902a,a6905a,a6909a,a6910a,a6911a,a6914a,a6918a,a6919a,a6920a,a6921a,a6922a,a6923a,a6924a,a6925a,a6926a,a6927a,a6928a,a6932a,a6933a,a6937a,a6938a,a6942a,a6943a,a6947a,a6948a,a6952a,a6953a,a6957a,a6958a,a6962a,a6963a,a6967a,a6968a,a6972a,a6973a,a6977a,a6978a,a6982a,a6983a,a6987a,a6988a,a6992a,a6993a,a6997a,a6998a,a7002a,a7003a,a7007a,a7008a,a7012a,a7013a,a7016a,a7019a,a7020a,a7024a,a7025a,a7028a,a7031a,a7032a,a7036a,a7037a,a7040a,a7043a,a7044a,a7048a,a7049a,a7052a,a7055a,a7056a,a7060a,a7061a,a7064a,a7067a,a7068a,a7072a,a7073a,a7076a,a7079a,a7080a,a7084a,a7085a,a7088a,a7091a,a7092a,a7096a,a7097a,a7100a,a7103a,a7104a,a7108a,a7109a,a7112a,a7115a,a7116a,a7120a,a7121a,a7124a,a7127a,a7128a,a7132a,a7133a,a7136a,a7139a,a7140a,a7144a,a7145a,a7148a,a7151a,a7152a,a7156a,a7157a,a7160a,a7163a,a7164a,a7168a,a7169a,a7172a,a7175a,a7176a,a7180a,a7181a,a7184a,a7187a,a7188a,a7192a,a7193a,a7196a,a7199a,a7200a,a7204a,a7205a,a7208a,a7211a,a7212a,a7216a,a7217a,a7220a,a7223a,a7224a,a7228a,a7229a,a7232a,a7235a,a7236a,a7240a,a7241a,a7244a,a7247a,a7248a,a7252a,a7253a,a7256a,a7259a,a7260a,a7264a,a7265a,a7268a,a7271a,a7272a,a7276a,a7277a,a7280a,a7283a,a7284a,a7288a,a7289a,a7292a,a7295a,a7296a,a7300a,a7301a,a7304a,a7307a,a7308a,a7312a,a7313a,a7316a,a7319a,a7320a,a7324a,a7325a,a7328a,a7331a,a7332a,a7336a,a7337a,a7340a,a7343a,a7344a,a7348a,a7349a,a7352a,a7355a,a7356a,a7360a,a7361a,a7364a,a7367a,a7368a,a7372a,a7373a,a7376a,a7379a,a7380a,a7384a,a7385a,a7388a,a7391a,a7392a,a7396a,a7397a,a7400a,a7403a,a7404a,a7408a,a7409a,a7412a,a7415a,a7416a,a7420a,a7421a,a7424a,a7427a,a7428a,a7432a,a7433a,a7436a,a7439a,a7440a,a7444a,a7445a,a7448a,a7451a,a7452a,a7456a,a7457a,a7460a,a7463a,a7464a,a7468a,a7469a,a7472a,a7475a,a7476a,a7480a,a7481a,a7484a,a7487a,a7488a,a7492a,a7493a,a7496a,a7499a,a7500a,a7504a,a7505a,a7508a,a7511a,a7512a,a7516a,a7517a,a7520a,a7523a,a7524a,a7528a,a7529a,a7532a,a7535a,a7536a,a7540a,a7541a,a7544a,a7547a,a7548a,a7552a,a7553a,a7556a,a7559a,a7560a,a7564a,a7565a,a7568a,a7571a,a7572a,a7576a,a7577a,a7580a,a7583a,a7584a,a7588a,a7589a,a7592a,a7595a,a7596a,a7600a,a7601a,a7604a,a7607a,a7608a,a7612a,a7613a,a7616a,a7619a,a7620a,a7624a,a7625a,a7628a,a7631a,a7632a,a7635a,a7638a,a7639a,a7642a,a7645a,a7646a,a7649a,a7652a,a7653a,a7656a,a7659a,a7660a,a7663a,a7666a,a7667a,a7670a,a7673a,a7674a,a7677a,a7680a,a7681a,a7684a,a7687a,a7688a,a7691a,a7694a,a7695a,a7698a,a7701a,a7702a,a7705a,a7708a,a7709a,a7712a,a7715a,a7716a,a7719a,a7722a,a7723a,a7726a,a7729a,a7730a,a7733a,a7736a,a7737a,a7740a,a7743a,a7744a,a7747a,a7750a,a7751a,a7754a,a7757a,a7758a,a7761a,a7764a,a7765a,a7768a,a7771a,a7772a,a7775a,a7778a,a7779a,a7782a,a7785a,a7786a,a7789a,a7792a,a7793a,a7796a,a7799a,a7800a,a7803a,a7806a,a7807a,a7810a,a7813a,a7814a,a7817a,a7820a,a7821a,a7824a,a7827a,a7828a,a7831a,a7834a,a7835a,a7838a,a7841a,a7842a,a7845a,a7848a,a7849a,a7852a,a7855a,a7856a,a7859a,a7862a,a7863a,a7866a,a7869a,a7870a,a7873a,a7876a,a7877a,a7880a,a7883a,a7884a,a7887a,a7890a,a7891a,a7894a,a7897a,a7898a,a7901a,a7904a,a7905a,a7908a,a7911a,a7912a,a7915a,a7918a,a7919a,a7922a,a7925a,a7926a,a7929a,a7932a,a7933a,a7936a,a7939a,a7940a,a7943a,a7946a,a7947a,a7950a,a7953a,a7954a,a7957a,a7960a,a7961a,a7964a,a7967a,a7968a,a7971a,a7974a,a7975a,a7978a,a7981a,a7982a,a7985a,a7988a,a7989a,a7992a,a7995a,a7996a,a7999a,a8002a,a8003a,a8006a,a8009a,a8010a,a8013a,a8016a,a8017a,a8020a,a8023a,a8024a,a8027a,a8030a,a8031a,a8034a,a8037a,a8038a,a8041a,a8044a,a8045a,a8048a,a8051a,a8052a,a8055a,a8058a,a8059a,a8062a,a8065a,a8066a,a8069a,a8072a,a8073a,a8076a,a8079a,a8080a,a8083a,a8086a,a8087a,a8090a,a8093a,a8094a,a8097a,a8100a,a8101a,a8104a,a8107a,a8108a,a8111a,a8114a,a8115a,a8118a,a8121a,a8122a,a8125a,a8128a,a8129a,a8132a,a8135a,a8136a,a8139a,a8142a,a8143a,a8146a,a8149a,a8150a,a8153a,a8156a,a8157a,a8160a,a8163a,a8164a,a8167a,a8170a,a8171a,a8174a,a8177a,a8178a,a8181a,a8184a,a8185a,a8188a,a8191a,a8192a,a8195a,a8198a,a8199a,a8202a,a8205a,a8206a,a8209a,a8212a,a8213a,a8216a,a8219a,a8220a,a8223a,a8226a,a8227a,a8230a,a8233a,a8234a,a8237a,a8240a,a8241a,a8244a,a8247a,a8248a,a8251a,a8254a,a8255a,a8258a,a8261a,a8262a,a8265a,a8268a,a8269a,a8272a,a8275a,a8276a,a8279a,a8282a,a8283a,a8286a,a8289a,a8290a,a8293a,a8296a,a8297a,a8300a,a8303a,a8304a,a8307a,a8310a,a8311a,a8314a,a8317a,a8318a,a8321a,a8324a,a8325a,a8328a,a8331a,a8332a,a8335a,a8338a,a8339a,a8342a,a8345a,a8346a,a8349a,a8352a,a8353a,a8356a,a8359a,a8360a,a8363a,a8366a,a8367a,a8370a,a8373a,a8374a,a8377a,a8380a,a8381a,a8384a,a8387a,a8388a,a8391a,a8394a,a8395a,a8398a,a8401a,a8402a,a8405a,a8408a,a8409a,a8412a,a8415a,a8416a,a8419a,a8422a,a8423a,a8426a,a8429a,a8430a,a8433a,a8436a,a8437a,a8440a,a8443a,a8444a,a8447a,a8450a,a8451a,a8454a,a8457a,a8458a,a8461a,a8464a,a8465a,a8468a,a8471a,a8472a,a8475a,a8478a,a8479a,a8482a,a8485a,a8486a,a8489a,a8492a,a8493a,a8496a,a8499a,a8500a,a8503a,a8506a,a8507a,a8510a,a8513a,a8514a,a8517a,a8520a,a8521a,a8524a,a8527a,a8528a,a8531a,a8534a,a8535a,a8538a,a8541a,a8542a,a8545a,a8548a,a8549a,a8552a,a8555a,a8556a,a8559a,a8562a,a8563a,a8566a,a8569a,a8570a,a8573a,a8576a,a8577a,a8580a,a8583a,a8584a,a8587a,a8590a,a8591a,a8594a,a8597a,a8598a,a8601a,a8604a,a8605a,a8608a,a8611a,a8612a,a8615a,a8618a,a8619a,a8622a,a8625a,a8626a,a8629a,a8632a,a8633a,a8636a,a8639a,a8640a,a8643a,a8646a,a8647a,a8650a,a8653a,a8654a,a8657a,a8660a,a8661a,a8664a,a8667a,a8668a,a8671a,a8674a,a8675a,a8678a,a8681a,a8682a,a8685a,a8688a,a8689a,a8692a,a8695a,a8696a,a8699a,a8702a,a8703a,a8706a,a8709a,a8710a,a8713a,a8716a,a8717a,a8720a,a8723a,a8724a,a8727a,a8730a,a8731a,a8734a,a8737a,a8738a,a8741a,a8744a,a8745a,a8748a,a8751a,a8752a,a8755a,a8758a,a8759a,a8762a,a8765a,a8766a,a8769a,a8772a,a8773a,a8776a,a8779a,a8780a,a8783a,a8786a,a8787a,a8790a,a8793a,a8794a,a8797a,a8800a,a8801a,a8804a,a8807a,a8808a,a8811a,a8814a,a8815a,a8818a,a8821a,a8822a,a8825a,a8828a,a8829a,a8832a,a8835a,a8836a,a8839a,a8842a,a8843a,a8846a,a8849a,a8850a,a8853a,a8856a,a8857a,a8860a,a8863a,a8864a,a8867a,a8870a,a8871a,a8874a,a8877a,a8878a,a8881a,a8884a,a8885a,a8888a,a8891a,a8892a,a8895a,a8898a,a8899a,a8902a,a8905a,a8906a,a8909a,a8912a,a8913a,a8916a,a8919a,a8920a,a8923a,a8926a,a8927a,a8930a,a8933a,a8934a,a8937a,a8940a,a8941a,a8944a,a8947a,a8948a,a8951a,a8954a,a8955a,a8958a,a8961a,a8962a,a8965a,a8968a,a8969a,a8972a,a8975a,a8976a,a8979a,a8982a,a8983a,a8986a,a8989a,a8990a,a8993a,a8996a,a8997a,a9000a,a9003a,a9004a,a9007a,a9010a,a9011a,a9014a,a9017a,a9018a,a9021a,a9024a,a9025a,a9028a,a9031a,a9032a,a9035a,a9038a,a9039a,a9042a,a9045a,a9046a,a9049a,a9052a,a9053a,a9056a,a9059a,a9060a,a9063a,a9066a,a9067a,a9070a,a9073a,a9074a,a9077a,a9080a,a9081a,a9084a,a9087a,a9088a,a9091a,a9094a,a9095a,a9098a,a9101a,a9102a,a9105a,a9108a,a9109a,a9112a,a9115a,a9116a,a9119a,a9122a,a9123a,a9126a,a9129a,a9130a,a9133a,a9136a,a9137a,a9140a,a9143a,a9144a,a9147a,a9150a,a9151a,a9154a,a9157a,a9158a,a9161a,a9164a,a9165a,a9168a,a9171a,a9172a,a9175a,a9178a,a9179a,a9182a,a9185a,a9186a,a9189a,a9192a,a9193a,a9196a,a9199a,a9200a,a9203a,a9206a,a9207a,a9210a,a9213a,a9214a,a9217a,a9220a,a9221a,a9224a,a9227a,a9228a,a9231a,a9234a,a9235a,a9238a,a9241a,a9242a,a9245a,a9248a,a9249a,a9252a,a9255a,a9256a,a9259a,a9262a,a9263a,a9266a,a9269a,a9270a,a9273a,a9276a,a9277a,a9280a,a9283a,a9284a,a9287a,a9290a,a9291a,a9294a,a9297a,a9298a,a9301a,a9304a,a9305a,a9308a,a9311a,a9312a,a9315a,a9318a,a9319a,a9322a,a9325a,a9326a,a9329a,a9332a,a9333a,a9336a,a9339a,a9340a,a9343a,a9346a,a9347a,a9350a,a9353a,a9354a,a9357a,a9360a,a9361a,a9364a,a9367a,a9368a,a9371a,a9374a,a9375a,a9378a,a9381a,a9382a,a9385a,a9388a,a9389a,a9392a,a9395a,a9396a,a9399a,a9402a,a9403a,a9406a,a9409a,a9410a,a9413a,a9416a,a9417a,a9420a,a9423a,a9424a,a9427a,a9430a,a9431a,a9434a,a9437a,a9438a,a9441a,a9444a,a9445a,a9448a,a9451a,a9452a,a9455a,a9458a,a9459a,a9462a,a9465a,a9466a,a9469a,a9472a,a9473a,a9476a,a9479a,a9480a,a9483a,a9486a,a9487a,a9490a,a9493a,a9494a,a9497a,a9500a,a9501a,a9504a,a9507a,a9508a,a9511a,a9514a,a9515a,a9518a,a9521a,a9522a,a9525a,a9528a,a9529a,a9532a,a9535a,a9536a,a9539a,a9542a,a9543a,a9546a,a9549a,a9550a,a9553a,a9556a,a9557a,a9560a,a9563a,a9564a,a9567a,a9570a,a9571a,a9574a,a9577a,a9578a,a9581a,a9584a,a9585a,a9588a,a9591a,a9592a,a9595a,a9598a,a9599a,a9602a,a9605a,a9606a,a9609a,a9612a,a9613a,a9616a,a9619a,a9620a,a9623a,a9626a,a9627a,a9630a,a9633a,a9634a,a9637a,a9640a,a9641a,a9644a,a9647a,a9648a,a9651a,a9654a,a9655a,a9658a,a9661a,a9662a,a9665a,a9668a,a9669a,a9672a,a9675a,a9676a,a9679a,a9682a,a9683a,a9686a,a9689a,a9690a,a9693a,a9696a,a9697a,a9700a,a9703a,a9704a,a9707a,a9710a,a9711a,a9714a,a9717a,a9718a,a9721a,a9724a,a9725a,a9728a,a9731a,a9732a,a9735a,a9738a,a9739a,a9742a,a9745a,a9746a,a9749a,a9752a,a9753a,a9756a,a9759a,a9760a,a9763a,a9766a,a9767a,a9770a,a9773a,a9774a,a9777a,a9780a,a9781a,a9784a,a9787a,a9788a,a9791a,a9794a,a9795a,a9798a,a9801a,a9802a,a9805a,a9808a,a9809a,a9812a,a9815a,a9816a,a9819a,a9822a,a9823a,a9826a,a9829a,a9830a,a9833a,a9836a,a9837a,a9840a,a9843a,a9844a,a9847a,a9850a,a9851a,a9854a,a9857a,a9858a,a9861a,a9864a,a9865a,a9868a,a9871a,a9872a,a9875a,a9878a,a9879a,a9882a,a9885a,a9886a,a9889a,a9892a,a9893a,a9896a,a9899a,a9900a,a9903a,a9906a,a9907a,a9910a,a9913a,a9914a,a9917a,a9920a,a9921a,a9924a,a9927a,a9928a,a9931a,a9934a,a9935a,a9938a,a9941a,a9942a,a9945a,a9948a,a9949a,a9952a,a9955a,a9956a,a9959a,a9962a,a9963a,a9966a,a9969a,a9970a,a9973a,a9976a,a9977a,a9980a,a9983a,a9984a,a9987a,a9990a,a9991a,a9994a,a9998a,a9999a,a10000a,a10003a,a10006a,a10007a,a10010a,a10014a,a10015a,a10016a,a10019a,a10022a,a10023a,a10026a,a10030a,a10031a,a10032a,a10035a,a10038a,a10039a,a10042a,a10046a,a10047a,a10048a,a10051a,a10054a,a10055a,a10058a,a10062a,a10063a,a10064a,a10067a,a10070a,a10071a,a10074a,a10078a,a10079a,a10080a,a10083a,a10086a,a10087a,a10090a,a10094a,a10095a,a10096a,a10099a,a10102a,a10103a,a10106a,a10110a,a10111a,a10112a,a10115a,a10118a,a10119a,a10122a,a10126a,a10127a,a10128a,a10131a,a10134a,a10135a,a10138a,a10142a,a10143a,a10144a,a10147a,a10150a,a10151a,a10154a,a10158a,a10159a,a10160a,a10163a,a10166a,a10167a,a10170a,a10174a,a10175a,a10176a,a10179a,a10182a,a10183a,a10186a,a10190a,a10191a,a10192a,a10195a,a10198a,a10199a,a10202a,a10206a,a10207a,a10208a,a10211a,a10214a,a10215a,a10218a,a10222a,a10223a,a10224a,a10227a,a10230a,a10231a,a10234a,a10238a,a10239a,a10240a,a10243a,a10246a,a10247a,a10250a,a10254a,a10255a,a10256a,a10259a,a10262a,a10263a,a10266a,a10270a,a10271a,a10272a,a10275a,a10278a,a10279a,a10282a,a10286a,a10287a,a10288a,a10291a,a10294a,a10295a,a10298a,a10302a,a10303a,a10304a,a10307a,a10310a,a10311a,a10314a,a10318a,a10319a,a10320a,a10323a,a10326a,a10327a,a10330a,a10334a,a10335a,a10336a,a10339a,a10342a,a10343a,a10346a,a10350a,a10351a,a10352a,a10355a,a10358a,a10359a,a10362a,a10366a,a10367a,a10368a,a10371a,a10374a,a10375a,a10378a,a10382a,a10383a,a10384a,a10387a,a10390a,a10391a,a10394a,a10398a,a10399a,a10400a,a10403a,a10406a,a10407a,a10410a,a10414a,a10415a,a10416a,a10419a,a10422a,a10423a,a10426a,a10430a,a10431a,a10432a,a10435a,a10438a,a10439a,a10442a,a10446a,a10447a,a10448a,a10451a,a10454a,a10455a,a10458a,a10462a,a10463a,a10464a,a10467a,a10470a,a10471a,a10474a,a10478a,a10479a,a10480a,a10483a,a10486a,a10487a,a10490a,a10494a,a10495a,a10496a,a10499a,a10502a,a10503a,a10506a,a10510a,a10511a,a10512a,a10515a,a10518a,a10519a,a10522a,a10526a,a10527a,a10528a,a10531a,a10534a,a10535a,a10538a,a10542a,a10543a,a10544a,a10547a,a10550a,a10551a,a10554a,a10558a,a10559a,a10560a,a10563a,a10566a,a10567a,a10570a,a10574a,a10575a,a10576a,a10579a,a10582a,a10583a,a10586a,a10590a,a10591a,a10592a,a10595a,a10598a,a10599a,a10602a,a10606a,a10607a,a10608a,a10611a,a10614a,a10615a,a10618a,a10622a,a10623a,a10624a,a10627a,a10630a,a10631a,a10634a,a10638a,a10639a,a10640a,a10643a,a10646a,a10647a,a10650a,a10654a,a10655a,a10656a,a10659a,a10662a,a10663a,a10666a,a10670a,a10671a,a10672a,a10675a,a10678a,a10679a,a10682a,a10686a,a10687a,a10688a,a10691a,a10694a,a10695a,a10698a,a10702a,a10703a,a10704a,a10707a,a10710a,a10711a,a10714a,a10718a,a10719a,a10720a,a10723a,a10726a,a10727a,a10730a,a10734a,a10735a,a10736a,a10739a,a10742a,a10743a,a10746a,a10750a,a10751a,a10752a,a10755a,a10758a,a10759a,a10762a,a10766a,a10767a,a10768a,a10771a,a10774a,a10775a,a10778a,a10782a,a10783a,a10784a,a10787a,a10790a,a10791a,a10794a,a10798a,a10799a,a10800a,a10803a,a10806a,a10807a,a10810a,a10814a,a10815a,a10816a,a10819a,a10822a,a10823a,a10826a,a10830a,a10831a,a10832a,a10835a,a10838a,a10839a,a10842a,a10846a,a10847a,a10848a,a10851a,a10854a,a10855a,a10858a,a10862a,a10863a,a10864a,a10867a,a10870a,a10871a,a10874a,a10878a,a10879a,a10880a,a10883a,a10886a,a10887a,a10890a,a10894a,a10895a,a10896a,a10899a,a10902a,a10903a,a10906a,a10910a,a10911a,a10912a,a10915a,a10918a,a10919a,a10922a,a10926a,a10927a,a10928a,a10931a,a10934a,a10935a,a10938a,a10942a,a10943a,a10944a,a10947a,a10950a,a10951a,a10954a,a10958a,a10959a,a10960a,a10963a,a10966a,a10967a,a10970a,a10974a,a10975a,a10976a,a10979a,a10982a,a10983a,a10986a,a10990a,a10991a,a10992a,a10995a,a10998a,a10999a,a11002a,a11006a,a11007a,a11008a,a11011a,a11014a,a11015a,a11018a,a11022a,a11023a,a11024a,a11027a,a11030a,a11031a,a11034a,a11038a,a11039a,a11040a,a11043a,a11046a,a11047a,a11050a,a11054a,a11055a,a11056a,a11059a,a11062a,a11063a,a11066a,a11070a,a11071a,a11072a,a11075a,a11078a,a11079a,a11082a,a11086a,a11087a,a11088a,a11091a,a11094a,a11095a,a11098a,a11102a,a11103a,a11104a,a11107a,a11110a,a11111a,a11114a,a11118a,a11119a,a11120a,a11123a,a11126a,a11127a,a11130a,a11134a,a11135a,a11136a,a11139a,a11142a,a11143a,a11146a,a11150a,a11151a,a11152a,a11155a,a11158a,a11159a,a11162a,a11166a,a11167a,a11168a,a11171a,a11174a,a11175a,a11178a,a11182a,a11183a,a11184a,a11187a,a11190a,a11191a,a11194a,a11198a,a11199a,a11200a,a11203a,a11206a,a11207a,a11210a,a11214a,a11215a,a11216a,a11219a,a11222a,a11223a,a11226a,a11230a,a11231a,a11232a,a11235a,a11238a,a11239a,a11242a,a11246a,a11247a,a11248a,a11251a,a11254a,a11255a,a11258a,a11262a,a11263a,a11264a,a11267a,a11270a,a11271a,a11274a,a11278a,a11279a,a11280a,a11283a,a11286a,a11287a,a11290a,a11294a,a11295a,a11296a,a11299a,a11302a,a11303a,a11306a,a11310a,a11311a,a11312a,a11315a,a11318a,a11319a,a11322a,a11326a,a11327a,a11328a,a11331a,a11334a,a11335a,a11338a,a11342a,a11343a,a11344a,a11347a,a11350a,a11351a,a11354a,a11358a,a11359a,a11360a,a11363a,a11366a,a11367a,a11370a,a11374a,a11375a,a11376a,a11379a,a11382a,a11383a,a11386a,a11390a,a11391a,a11392a,a11395a,a11398a,a11399a,a11402a,a11406a,a11407a,a11408a,a11411a,a11414a,a11415a,a11418a,a11422a,a11423a,a11424a,a11427a,a11430a,a11431a,a11434a,a11438a,a11439a,a11440a,a11443a,a11446a,a11447a,a11450a,a11454a,a11455a,a11456a,a11459a,a11462a,a11463a,a11466a,a11470a,a11471a,a11472a,a11475a,a11478a,a11479a,a11482a,a11486a,a11487a,a11488a,a11491a,a11494a,a11495a,a11498a,a11502a,a11503a,a11504a,a11507a,a11510a,a11511a,a11514a,a11518a,a11519a,a11520a,a11523a,a11526a,a11527a,a11530a,a11534a,a11535a,a11536a,a11539a,a11542a,a11543a,a11546a,a11550a,a11551a,a11552a,a11555a,a11558a,a11559a,a11562a,a11566a,a11567a,a11568a,a11571a,a11574a,a11575a,a11578a,a11582a,a11583a,a11584a,a11587a,a11590a,a11591a,a11594a,a11598a,a11599a,a11600a,a11603a,a11606a,a11607a,a11610a,a11614a,a11615a,a11616a,a11619a,a11622a,a11623a,a11626a,a11630a,a11631a,a11632a,a11635a,a11638a,a11639a,a11642a,a11646a,a11647a,a11648a,a11651a,a11654a,a11655a,a11658a,a11662a,a11663a,a11664a,a11667a,a11670a,a11671a,a11674a,a11678a,a11679a,a11680a,a11683a,a11686a,a11687a,a11690a,a11694a,a11695a,a11696a,a11699a,a11702a,a11703a,a11706a,a11710a,a11711a,a11712a,a11715a,a11718a,a11719a,a11722a,a11726a,a11727a,a11728a,a11731a,a11734a,a11735a,a11738a,a11742a,a11743a,a11744a,a11747a,a11750a,a11751a,a11754a,a11758a,a11759a,a11760a,a11763a,a11766a,a11767a,a11770a,a11774a,a11775a,a11776a,a11779a,a11782a,a11783a,a11786a,a11790a,a11791a,a11792a,a11795a,a11798a,a11799a,a11802a,a11806a,a11807a,a11808a,a11811a,a11814a,a11815a,a11818a,a11822a,a11823a,a11824a,a11827a,a11830a,a11831a,a11834a,a11838a,a11839a,a11840a,a11843a,a11846a,a11847a,a11850a,a11854a,a11855a,a11856a,a11859a,a11862a,a11863a,a11866a,a11870a,a11871a,a11872a,a11875a,a11878a,a11879a,a11882a,a11886a,a11887a,a11888a,a11891a,a11894a,a11895a,a11898a,a11902a,a11903a,a11904a,a11907a,a11910a,a11911a,a11914a,a11918a,a11919a,a11920a,a11923a,a11926a,a11927a,a11930a,a11934a,a11935a,a11936a,a11939a,a11942a,a11943a,a11946a,a11950a,a11951a,a11952a,a11955a,a11958a,a11959a,a11962a,a11966a,a11967a,a11968a,a11971a,a11974a,a11975a,a11978a,a11982a,a11983a,a11984a,a11987a,a11990a,a11991a,a11994a,a11998a,a11999a,a12000a,a12003a,a12006a,a12007a,a12010a,a12014a,a12015a,a12016a,a12019a,a12022a,a12023a,a12026a,a12030a,a12031a,a12032a,a12035a,a12038a,a12039a,a12042a,a12046a,a12047a,a12048a,a12051a,a12054a,a12055a,a12058a,a12062a,a12063a,a12064a,a12067a,a12070a,a12071a,a12074a,a12078a,a12079a,a12080a,a12083a,a12086a,a12087a,a12090a,a12094a,a12095a,a12096a,a12099a,a12102a,a12103a,a12106a,a12110a,a12111a,a12112a,a12115a,a12118a,a12119a,a12122a,a12126a,a12127a,a12128a,a12131a,a12134a,a12135a,a12138a,a12142a,a12143a,a12144a,a12147a,a12150a,a12151a,a12154a,a12158a,a12159a,a12160a,a12163a,a12166a,a12167a,a12170a,a12174a,a12175a,a12176a,a12179a,a12182a,a12183a,a12186a,a12190a,a12191a,a12192a,a12195a,a12198a,a12199a,a12202a,a12206a,a12207a,a12208a,a12211a,a12214a,a12215a,a12218a,a12222a,a12223a,a12224a,a12227a,a12230a,a12231a,a12234a,a12238a,a12239a,a12240a,a12243a,a12246a,a12247a,a12250a,a12254a,a12255a,a12256a,a12259a,a12262a,a12263a,a12266a,a12270a,a12271a,a12272a,a12275a,a12278a,a12279a,a12282a,a12286a,a12287a,a12288a,a12291a,a12294a,a12295a,a12298a,a12302a,a12303a,a12304a,a12307a,a12310a,a12311a,a12314a,a12318a,a12319a,a12320a,a12323a,a12326a,a12327a,a12330a,a12334a,a12335a,a12336a,a12339a,a12342a,a12343a,a12346a,a12350a,a12351a,a12352a,a12355a,a12358a,a12359a,a12362a,a12366a,a12367a,a12368a,a12371a,a12374a,a12375a,a12378a,a12382a,a12383a,a12384a,a12387a,a12390a,a12391a,a12394a,a12398a,a12399a,a12400a,a12403a,a12406a,a12407a,a12410a,a12414a,a12415a,a12416a,a12419a,a12422a,a12423a,a12426a,a12430a,a12431a,a12432a,a12435a,a12438a,a12439a,a12442a,a12446a,a12447a,a12448a,a12451a,a12454a,a12455a,a12458a,a12462a,a12463a,a12464a,a12467a,a12470a,a12471a,a12474a,a12478a,a12479a,a12480a,a12483a,a12486a,a12487a,a12490a,a12494a,a12495a,a12496a,a12499a,a12502a,a12503a,a12506a,a12510a,a12511a,a12512a,a12515a,a12518a,a12519a,a12522a,a12526a,a12527a,a12528a,a12531a,a12534a,a12535a,a12538a,a12542a,a12543a,a12544a,a12547a,a12550a,a12551a,a12554a,a12558a,a12559a,a12560a,a12563a,a12566a,a12567a,a12570a,a12574a,a12575a,a12576a,a12579a,a12582a,a12583a,a12586a,a12590a,a12591a,a12592a,a12595a,a12598a,a12599a,a12602a,a12606a,a12607a,a12608a,a12611a,a12614a,a12615a,a12618a,a12622a,a12623a,a12624a,a12627a,a12630a,a12631a,a12634a,a12638a,a12639a,a12640a,a12643a,a12646a,a12647a,a12650a,a12654a,a12655a,a12656a,a12659a,a12662a,a12663a,a12666a,a12670a,a12671a,a12672a,a12675a,a12678a,a12679a,a12682a,a12686a,a12687a,a12688a,a12691a,a12694a,a12695a,a12698a,a12702a,a12703a,a12704a,a12707a,a12710a,a12711a,a12714a,a12718a,a12719a,a12720a,a12723a,a12726a,a12727a,a12730a,a12734a,a12735a,a12736a,a12739a,a12742a,a12743a,a12746a,a12750a,a12751a,a12752a,a12755a,a12758a,a12759a,a12762a,a12766a,a12767a,a12768a,a12771a,a12774a,a12775a,a12778a,a12782a,a12783a,a12784a,a12787a,a12790a,a12791a,a12794a,a12798a,a12799a,a12800a,a12803a,a12806a,a12807a,a12810a,a12814a,a12815a,a12816a,a12819a,a12822a,a12823a,a12826a,a12830a,a12831a,a12832a,a12835a,a12838a,a12839a,a12842a,a12846a,a12847a,a12848a,a12851a,a12854a,a12855a,a12858a,a12862a,a12863a,a12864a,a12867a,a12870a,a12871a,a12874a,a12878a,a12879a,a12880a,a12883a,a12886a,a12887a,a12890a,a12894a,a12895a,a12896a,a12899a,a12902a,a12903a,a12906a,a12910a,a12911a,a12912a,a12915a,a12918a,a12919a,a12922a,a12926a,a12927a,a12928a,a12931a,a12934a,a12935a,a12938a,a12942a,a12943a,a12944a,a12947a,a12950a,a12951a,a12954a,a12958a,a12959a,a12960a,a12963a,a12966a,a12967a,a12970a,a12974a,a12975a,a12976a,a12979a,a12982a,a12983a,a12986a,a12990a,a12991a,a12992a,a12995a,a12998a,a12999a,a13002a,a13006a,a13007a,a13008a,a13011a,a13014a,a13015a,a13018a,a13022a,a13023a,a13024a,a13027a,a13030a,a13031a,a13034a,a13038a,a13039a,a13040a,a13043a,a13046a,a13047a,a13050a,a13054a,a13055a,a13056a,a13059a,a13062a,a13063a,a13066a,a13070a,a13071a,a13072a,a13075a,a13078a,a13079a,a13082a,a13086a,a13087a,a13088a,a13091a,a13094a,a13095a,a13098a,a13102a,a13103a,a13104a,a13107a,a13110a,a13111a,a13114a,a13118a,a13119a,a13120a,a13123a,a13126a,a13127a,a13130a,a13134a,a13135a,a13136a,a13139a,a13142a,a13143a,a13146a,a13150a,a13151a,a13152a,a13155a,a13158a,a13159a,a13162a,a13166a,a13167a,a13168a,a13171a,a13174a,a13175a,a13178a,a13182a,a13183a,a13184a,a13187a,a13190a,a13191a,a13194a,a13198a,a13199a,a13200a,a13203a,a13206a,a13207a,a13210a,a13214a,a13215a,a13216a,a13219a,a13222a,a13223a,a13226a,a13230a,a13231a,a13232a,a13235a,a13238a,a13239a,a13242a,a13246a,a13247a,a13248a,a13251a,a13254a,a13255a,a13258a,a13262a,a13263a,a13264a,a13267a,a13270a,a13271a,a13274a,a13278a,a13279a,a13280a,a13283a,a13286a,a13287a,a13290a,a13294a,a13295a,a13296a,a13299a,a13302a,a13303a,a13306a,a13310a,a13311a,a13312a,a13315a,a13318a,a13319a,a13322a,a13326a,a13327a,a13328a,a13331a,a13334a,a13335a,a13338a,a13342a,a13343a,a13344a,a13347a,a13350a,a13351a,a13354a,a13358a,a13359a,a13360a,a13363a,a13366a,a13367a,a13370a,a13374a,a13375a,a13376a,a13379a,a13382a,a13383a,a13386a,a13390a,a13391a,a13392a,a13395a,a13398a,a13399a,a13402a,a13406a,a13407a,a13408a,a13411a,a13414a,a13415a,a13418a,a13422a,a13423a,a13424a,a13427a,a13430a,a13431a,a13434a,a13438a,a13439a,a13440a,a13443a,a13446a,a13447a,a13450a,a13454a,a13455a,a13456a,a13459a,a13462a,a13463a,a13466a,a13470a,a13471a,a13472a,a13475a,a13478a,a13479a,a13482a,a13486a,a13487a,a13488a,a13491a,a13494a,a13495a,a13498a,a13502a,a13503a,a13504a,a13507a,a13510a,a13511a,a13514a,a13518a,a13519a,a13520a,a13523a,a13526a,a13527a,a13530a,a13534a,a13535a,a13536a,a13539a,a13542a,a13543a,a13546a,a13550a,a13551a,a13552a,a13555a,a13558a,a13559a,a13562a,a13566a,a13567a,a13568a,a13571a,a13574a,a13575a,a13578a,a13582a,a13583a,a13584a,a13587a,a13590a,a13591a,a13594a,a13598a,a13599a,a13600a,a13603a,a13606a,a13607a,a13610a,a13614a,a13615a,a13616a,a13619a,a13622a,a13623a,a13626a,a13630a,a13631a,a13632a,a13635a,a13638a,a13639a,a13642a,a13646a,a13647a,a13648a,a13651a,a13654a,a13655a,a13658a,a13662a,a13663a,a13664a,a13667a,a13670a,a13671a,a13674a,a13678a,a13679a,a13680a,a13683a,a13686a,a13687a,a13690a,a13694a,a13695a,a13696a,a13699a,a13702a,a13703a,a13706a,a13710a,a13711a,a13712a,a13715a,a13718a,a13719a,a13722a,a13726a,a13727a,a13728a,a13731a,a13734a,a13735a,a13738a,a13742a,a13743a,a13744a,a13747a,a13750a,a13751a,a13754a,a13758a,a13759a,a13760a,a13763a,a13766a,a13767a,a13770a,a13774a,a13775a,a13776a,a13779a,a13782a,a13783a,a13786a,a13790a,a13791a,a13792a,a13795a,a13798a,a13799a,a13802a,a13806a,a13807a,a13808a,a13811a,a13814a,a13815a,a13818a,a13822a,a13823a,a13824a,a13827a,a13830a,a13831a,a13834a,a13838a,a13839a,a13840a,a13843a,a13846a,a13847a,a13850a,a13854a,a13855a,a13856a,a13859a,a13862a,a13863a,a13866a,a13870a,a13871a,a13872a,a13875a,a13878a,a13879a,a13882a,a13886a,a13887a,a13888a,a13891a,a13894a,a13895a,a13898a,a13902a,a13903a,a13904a,a13907a,a13910a,a13911a,a13914a,a13918a,a13919a,a13920a,a13923a,a13926a,a13927a,a13930a,a13934a,a13935a,a13936a,a13939a,a13942a,a13943a,a13946a,a13950a,a13951a,a13952a,a13955a,a13958a,a13959a,a13962a,a13966a,a13967a,a13968a,a13971a,a13974a,a13975a,a13978a,a13982a,a13983a,a13984a,a13987a,a13990a,a13991a,a13994a,a13998a,a13999a,a14000a,a14003a,a14006a,a14007a,a14010a,a14014a,a14015a,a14016a,a14019a,a14022a,a14023a,a14026a,a14030a,a14031a,a14032a,a14035a,a14038a,a14039a,a14042a,a14046a,a14047a,a14048a,a14051a,a14054a,a14055a,a14058a,a14062a,a14063a,a14064a,a14067a,a14070a,a14071a,a14074a,a14078a,a14079a,a14080a,a14083a,a14086a,a14087a,a14090a,a14094a,a14095a,a14096a,a14099a,a14102a,a14103a,a14106a,a14110a,a14111a,a14112a,a14115a,a14118a,a14119a,a14122a,a14126a,a14127a,a14128a,a14131a,a14134a,a14135a,a14138a,a14142a,a14143a,a14144a,a14147a,a14150a,a14151a,a14154a,a14158a,a14159a,a14160a,a14163a,a14166a,a14167a,a14170a,a14174a,a14175a,a14176a,a14179a,a14182a,a14183a,a14186a,a14190a,a14191a,a14192a,a14195a,a14198a,a14199a,a14202a,a14206a,a14207a,a14208a,a14211a,a14214a,a14215a,a14218a,a14222a,a14223a,a14224a,a14227a,a14230a,a14231a,a14234a,a14238a,a14239a,a14240a,a14243a,a14246a,a14247a,a14250a,a14254a,a14255a,a14256a,a14259a,a14262a,a14263a,a14266a,a14270a,a14271a,a14272a,a14275a,a14278a,a14279a,a14282a,a14286a,a14287a,a14288a,a14291a,a14294a,a14295a,a14298a,a14302a,a14303a,a14304a,a14307a,a14310a,a14311a,a14314a,a14318a,a14319a,a14320a,a14323a,a14326a,a14327a,a14330a,a14334a,a14335a,a14336a,a14339a,a14342a,a14343a,a14346a,a14350a,a14351a,a14352a,a14355a,a14358a,a14359a,a14362a,a14366a,a14367a,a14368a,a14371a,a14374a,a14375a,a14378a,a14382a,a14383a,a14384a,a14387a,a14390a,a14391a,a14394a,a14398a,a14399a,a14400a,a14403a,a14406a,a14407a,a14410a,a14414a,a14415a,a14416a,a14419a,a14422a,a14423a,a14426a,a14430a,a14431a,a14432a,a14435a,a14438a,a14439a,a14442a,a14446a,a14447a,a14448a,a14451a,a14454a,a14455a,a14458a,a14462a,a14463a,a14464a,a14467a,a14470a,a14471a,a14474a,a14478a,a14479a,a14480a,a14483a,a14486a,a14487a,a14490a,a14494a,a14495a,a14496a,a14499a,a14502a,a14503a,a14506a,a14510a,a14511a,a14512a,a14515a,a14518a,a14519a,a14522a,a14526a,a14527a,a14528a,a14531a,a14534a,a14535a,a14538a,a14542a,a14543a,a14544a,a14547a,a14550a,a14551a,a14554a,a14558a,a14559a,a14560a,a14563a,a14566a,a14567a,a14570a,a14574a,a14575a,a14576a,a14579a,a14582a,a14583a,a14586a,a14590a,a14591a,a14592a,a14595a,a14598a,a14599a,a14602a,a14606a,a14607a,a14608a,a14611a,a14614a,a14615a,a14618a,a14622a,a14623a,a14624a,a14627a,a14630a,a14631a,a14634a,a14638a,a14639a,a14640a,a14643a,a14646a,a14647a,a14650a,a14654a,a14655a,a14656a,a14659a,a14662a,a14663a,a14666a,a14670a,a14671a,a14672a,a14675a,a14678a,a14679a,a14682a,a14686a,a14687a,a14688a,a14691a,a14694a,a14695a,a14698a,a14702a,a14703a,a14704a,a14707a,a14710a,a14711a,a14714a,a14718a,a14719a,a14720a,a14723a,a14726a,a14727a,a14730a,a14734a,a14735a,a14736a,a14739a,a14742a,a14743a,a14746a,a14750a,a14751a,a14752a,a14755a,a14758a,a14759a,a14762a,a14766a,a14767a,a14768a,a14771a,a14774a,a14775a,a14778a,a14782a,a14783a,a14784a,a14787a,a14790a,a14791a,a14794a,a14798a,a14799a,a14800a,a14803a,a14806a,a14807a,a14810a,a14814a,a14815a,a14816a,a14819a,a14822a,a14823a,a14826a,a14830a,a14831a,a14832a,a14835a,a14838a,a14839a,a14842a,a14846a,a14847a,a14848a,a14851a,a14854a,a14855a,a14858a,a14862a,a14863a,a14864a,a14867a,a14870a,a14871a,a14874a,a14878a,a14879a,a14880a,a14883a,a14886a,a14887a,a14890a,a14894a,a14895a,a14896a,a14899a,a14902a,a14903a,a14906a,a14910a,a14911a,a14912a,a14915a,a14918a,a14919a,a14922a,a14926a,a14927a,a14928a,a14931a,a14934a,a14935a,a14938a,a14942a,a14943a,a14944a,a14947a,a14950a,a14951a,a14954a,a14958a,a14959a,a14960a,a14963a,a14966a,a14967a,a14970a,a14974a,a14975a,a14976a,a14979a,a14982a,a14983a,a14986a,a14990a,a14991a,a14992a,a14995a,a14998a,a14999a,a15002a,a15006a,a15007a,a15008a,a15011a,a15014a,a15015a,a15018a,a15022a,a15023a,a15024a,a15027a,a15030a,a15031a,a15034a,a15038a,a15039a,a15040a,a15043a,a15046a,a15047a,a15050a,a15054a,a15055a,a15056a,a15059a,a15062a,a15063a,a15066a,a15070a,a15071a,a15072a,a15075a,a15078a,a15079a,a15082a,a15086a,a15087a,a15088a,a15091a,a15094a,a15095a,a15098a,a15102a,a15103a,a15104a,a15107a,a15110a,a15111a,a15114a,a15118a,a15119a,a15120a,a15123a,a15126a,a15127a,a15130a,a15134a,a15135a,a15136a,a15139a,a15142a,a15143a,a15146a,a15150a,a15151a,a15152a,a15155a,a15158a,a15159a,a15162a,a15166a,a15167a,a15168a,a15171a,a15174a,a15175a,a15178a,a15182a,a15183a,a15184a,a15187a,a15190a,a15191a,a15194a,a15198a,a15199a,a15200a,a15203a,a15206a,a15207a,a15210a,a15214a,a15215a,a15216a,a15219a,a15222a,a15223a,a15226a,a15230a,a15231a,a15232a,a15235a,a15239a,a15240a,a15241a,a15244a,a15248a,a15249a,a15250a,a15253a,a15257a,a15258a,a15259a,a15262a,a15266a,a15267a,a15268a,a15271a,a15275a,a15276a,a15277a,a15280a,a15284a,a15285a,a15286a,a15289a,a15293a,a15294a,a15295a,a15298a,a15302a,a15303a,a15304a,a15307a,a15311a,a15312a,a15313a,a15316a,a15320a,a15321a,a15322a,a15325a,a15329a,a15330a,a15331a,a15334a,a15338a,a15339a,a15340a,a15343a,a15347a,a15348a,a15349a,a15352a,a15356a,a15357a,a15358a,a15361a,a15365a,a15366a,a15367a,a15370a,a15374a,a15375a,a15376a,a15379a,a15383a,a15384a,a15385a,a15388a,a15392a,a15393a,a15394a,a15397a,a15401a,a15402a,a15403a,a15406a,a15410a,a15411a,a15412a,a15415a,a15419a,a15420a,a15421a,a15424a,a15428a,a15429a,a15430a,a15433a,a15437a,a15438a,a15439a,a15442a,a15446a,a15447a,a15448a,a15451a,a15455a,a15456a,a15457a,a15460a,a15464a,a15465a,a15466a,a15469a,a15473a,a15474a,a15475a,a15478a,a15482a,a15483a,a15484a,a15487a,a15491a,a15492a,a15493a,a15496a,a15500a,a15501a,a15502a,a15505a,a15509a,a15510a,a15511a,a15514a,a15518a,a15519a,a15520a,a15523a,a15527a,a15528a,a15529a,a15532a,a15536a,a15537a,a15538a,a15541a,a15545a,a15546a,a15547a,a15550a,a15554a,a15555a,a15556a,a15559a,a15563a,a15564a,a15565a,a15568a,a15572a,a15573a,a15574a,a15577a,a15581a,a15582a,a15583a,a15586a,a15590a,a15591a,a15592a,a15595a,a15599a,a15600a,a15601a,a15604a,a15608a,a15609a,a15610a,a15613a,a15617a,a15618a,a15619a,a15622a,a15626a,a15627a,a15628a,a15631a,a15635a,a15636a,a15637a,a15640a,a15644a,a15645a,a15646a,a15649a,a15653a,a15654a,a15655a,a15658a,a15662a,a15663a,a15664a,a15667a,a15671a,a15672a,a15673a,a15676a,a15680a,a15681a,a15682a,a15685a,a15689a,a15690a,a15691a,a15694a,a15698a,a15699a,a15700a,a15703a,a15707a,a15708a,a15709a,a15712a,a15716a,a15717a,a15718a,a15721a,a15725a,a15726a,a15727a,a15730a,a15734a,a15735a,a15736a,a15739a,a15743a,a15744a,a15745a,a15748a,a15752a,a15753a,a15754a,a15757a,a15761a,a15762a,a15763a,a15766a,a15770a,a15771a,a15772a,a15775a,a15779a,a15780a,a15781a,a15784a,a15788a,a15789a,a15790a,a15793a,a15797a,a15798a,a15799a,a15802a,a15806a,a15807a,a15808a,a15811a,a15815a,a15816a,a15817a,a15820a,a15824a,a15825a,a15826a,a15829a,a15833a,a15834a,a15835a,a15838a,a15842a,a15843a,a15844a,a15847a,a15851a,a15852a,a15853a,a15856a,a15860a,a15861a,a15862a,a15865a,a15869a,a15870a,a15871a,a15874a,a15878a,a15879a,a15880a,a15883a,a15887a,a15888a,a15889a,a15892a,a15896a,a15897a,a15898a,a15901a,a15905a,a15906a,a15907a,a15910a,a15914a,a15915a,a15916a,a15919a,a15923a,a15924a,a15925a,a15928a,a15932a,a15933a,a15934a,a15937a,a15941a,a15942a,a15943a,a15946a,a15950a,a15951a,a15952a,a15955a,a15959a,a15960a,a15961a,a15964a,a15968a,a15969a,a15970a,a15973a,a15977a,a15978a,a15979a,a15982a,a15986a,a15987a,a15988a,a15991a,a15995a,a15996a,a15997a,a16000a,a16004a,a16005a,a16006a,a16009a,a16013a,a16014a,a16015a,a16018a,a16022a,a16023a,a16024a,a16027a,a16031a,a16032a,a16033a,a16036a,a16040a,a16041a,a16042a,a16045a,a16049a,a16050a,a16051a,a16054a,a16058a,a16059a,a16060a,a16063a,a16067a,a16068a,a16069a,a16072a,a16076a,a16077a,a16078a,a16081a,a16085a,a16086a,a16087a,a16090a,a16094a,a16095a,a16096a,a16099a,a16103a,a16104a,a16105a,a16108a,a16112a,a16113a,a16114a,a16117a,a16121a,a16122a,a16123a,a16126a,a16130a,a16131a,a16132a,a16135a,a16139a,a16140a,a16141a,a16144a,a16148a,a16149a,a16150a,a16153a,a16157a,a16158a,a16159a,a16162a,a16166a,a16167a,a16168a,a16171a,a16175a,a16176a,a16177a,a16180a,a16184a,a16185a,a16186a,a16189a,a16193a,a16194a,a16195a,a16198a,a16202a,a16203a,a16204a,a16207a,a16211a,a16212a,a16213a,a16216a,a16220a,a16221a,a16222a,a16225a,a16229a,a16230a,a16231a,a16234a,a16238a,a16239a,a16240a,a16243a,a16247a,a16248a,a16249a,a16252a,a16256a,a16257a,a16258a,a16261a,a16265a,a16266a,a16267a,a16270a,a16274a,a16275a,a16276a,a16279a,a16283a,a16284a,a16285a,a16288a,a16292a,a16293a,a16294a,a16297a,a16301a,a16302a,a16303a,a16306a,a16310a,a16311a,a16312a,a16315a,a16319a,a16320a,a16321a,a16324a,a16328a,a16329a,a16330a,a16333a,a16337a,a16338a,a16339a,a16342a,a16346a,a16347a,a16348a,a16351a,a16355a,a16356a,a16357a,a16360a,a16364a,a16365a,a16366a,a16369a,a16373a,a16374a,a16375a,a16378a,a16382a,a16383a,a16384a,a16387a,a16391a,a16392a,a16393a,a16396a,a16400a,a16401a,a16402a,a16405a,a16409a,a16410a,a16411a,a16414a,a16418a,a16419a,a16420a,a16423a,a16427a,a16428a,a16429a,a16432a,a16436a,a16437a,a16438a,a16441a,a16445a,a16446a,a16447a,a16450a,a16454a,a16455a,a16456a,a16459a,a16463a,a16464a,a16465a,a16468a,a16472a,a16473a,a16474a,a16477a,a16481a,a16482a,a16483a,a16486a,a16490a,a16491a,a16492a,a16495a,a16499a,a16500a,a16501a,a16504a,a16508a,a16509a,a16510a,a16513a,a16517a,a16518a,a16519a,a16522a,a16526a,a16527a,a16528a,a16531a,a16535a,a16536a,a16537a,a16540a,a16544a,a16545a,a16546a,a16549a,a16553a,a16554a,a16555a,a16558a,a16562a,a16563a,a16564a,a16567a,a16571a,a16572a,a16573a,a16576a,a16580a,a16581a,a16582a,a16585a,a16589a,a16590a,a16591a,a16594a,a16598a,a16599a,a16600a,a16603a,a16607a,a16608a,a16609a,a16612a,a16616a,a16617a,a16618a,a16621a,a16625a,a16626a,a16627a,a16630a,a16634a,a16635a,a16636a,a16639a,a16643a,a16644a,a16645a,a16648a,a16652a,a16653a,a16654a,a16657a,a16661a,a16662a,a16663a,a16666a,a16670a,a16671a,a16672a,a16675a,a16679a,a16680a,a16681a,a16684a,a16688a,a16689a,a16690a,a16693a,a16697a,a16698a,a16699a,a16702a,a16706a,a16707a,a16708a,a16711a,a16715a,a16716a,a16717a,a16720a,a16724a,a16725a,a16726a,a16729a,a16733a,a16734a,a16735a,a16738a,a16742a,a16743a,a16744a,a16747a,a16751a,a16752a,a16753a,a16756a,a16760a,a16761a,a16762a,a16765a,a16769a,a16770a,a16771a,a16774a,a16778a,a16779a,a16780a,a16783a,a16787a,a16788a,a16789a,a16792a,a16796a,a16797a,a16798a,a16801a,a16805a,a16806a,a16807a,a16810a,a16814a,a16815a,a16816a,a16819a,a16823a,a16824a,a16825a,a16828a,a16832a,a16833a,a16834a,a16837a,a16841a,a16842a,a16843a,a16846a,a16850a,a16851a,a16852a,a16855a,a16859a,a16860a,a16861a,a16864a,a16868a,a16869a,a16870a,a16873a,a16877a,a16878a,a16879a,a16882a,a16886a,a16887a,a16888a,a16891a,a16895a,a16896a,a16897a,a16900a,a16904a,a16905a,a16906a,a16909a,a16913a,a16914a,a16915a,a16918a,a16922a,a16923a,a16924a,a16927a,a16931a,a16932a,a16933a,a16936a,a16940a,a16941a,a16942a,a16945a,a16949a,a16950a,a16951a,a16954a,a16958a,a16959a,a16960a,a16963a,a16967a,a16968a,a16969a,a16972a,a16976a,a16977a,a16978a,a16981a,a16985a,a16986a,a16987a,a16990a,a16994a,a16995a,a16996a,a16999a,a17003a,a17004a,a17005a,a17008a,a17012a,a17013a,a17014a,a17017a,a17021a,a17022a,a17023a,a17026a,a17030a,a17031a,a17032a,a17035a,a17039a,a17040a,a17041a,a17044a,a17048a,a17049a,a17050a,a17053a,a17057a,a17058a,a17059a,a17062a,a17066a,a17067a,a17068a,a17071a,a17075a,a17076a,a17077a,a17080a,a17084a,a17085a,a17086a,a17089a,a17093a,a17094a,a17095a,a17098a,a17102a,a17103a,a17104a,a17107a,a17111a,a17112a,a17113a,a17116a,a17120a,a17121a,a17122a,a17125a,a17129a,a17130a,a17131a,a17134a,a17138a,a17139a,a17140a,a17143a,a17147a,a17148a,a17149a,a17152a,a17156a,a17157a,a17158a,a17161a,a17165a,a17166a,a17167a,a17170a,a17174a,a17175a,a17176a,a17179a,a17183a,a17184a,a17185a,a17188a,a17192a,a17193a,a17194a,a17197a,a17201a,a17202a,a17203a,a17206a,a17210a,a17211a,a17212a,a17215a,a17219a,a17220a,a17221a,a17224a,a17228a,a17229a,a17230a,a17233a,a17237a,a17238a,a17239a,a17242a,a17246a,a17247a,a17248a,a17251a,a17255a,a17256a,a17257a,a17260a,a17264a,a17265a,a17266a,a17269a,a17273a,a17274a,a17275a,a17278a,a17282a,a17283a,a17284a,a17287a,a17291a,a17292a,a17293a,a17296a,a17300a,a17301a,a17302a,a17305a,a17309a,a17310a,a17311a,a17314a,a17318a,a17319a,a17320a,a17323a,a17327a,a17328a,a17329a,a17332a,a17336a,a17337a,a17338a,a17341a,a17345a,a17346a,a17347a,a17350a,a17354a,a17355a,a17356a,a17359a,a17363a,a17364a,a17365a,a17368a,a17372a,a17373a,a17374a,a17377a,a17381a,a17382a,a17383a,a17386a,a17390a,a17391a,a17392a,a17395a,a17399a,a17400a,a17401a,a17404a,a17408a,a17409a,a17410a,a17413a,a17417a,a17418a,a17419a,a17422a,a17426a,a17427a,a17428a,a17431a,a17435a,a17436a,a17437a,a17440a,a17444a,a17445a,a17446a,a17449a,a17453a,a17454a,a17455a,a17458a,a17462a,a17463a,a17464a,a17467a,a17471a,a17472a,a17473a,a17476a,a17480a,a17481a,a17482a,a17485a,a17489a,a17490a,a17491a,a17494a,a17498a,a17499a,a17500a,a17503a,a17507a,a17508a,a17509a,a17512a,a17516a,a17517a,a17518a,a17521a,a17525a,a17526a,a17527a,a17530a,a17534a,a17535a,a17536a,a17539a,a17543a,a17544a,a17545a,a17548a,a17552a,a17553a,a17554a,a17557a,a17561a,a17562a,a17563a,a17566a,a17570a,a17571a,a17572a,a17575a,a17579a,a17580a,a17581a,a17584a,a17588a,a17589a,a17590a,a17593a,a17597a,a17598a,a17599a,a17602a,a17606a,a17607a,a17608a,a17611a,a17615a,a17616a,a17617a,a17620a,a17624a,a17625a,a17626a,a17629a,a17633a,a17634a,a17635a,a17638a,a17642a,a17643a,a17644a,a17647a,a17651a,a17652a,a17653a,a17656a,a17660a,a17661a,a17662a,a17665a,a17669a,a17670a,a17671a,a17674a,a17678a,a17679a,a17680a,a17683a,a17687a,a17688a,a17689a,a17692a,a17696a,a17697a,a17698a,a17701a,a17705a,a17706a,a17707a,a17710a,a17714a,a17715a,a17716a,a17719a,a17723a,a17724a,a17725a,a17728a,a17732a,a17733a,a17734a,a17737a,a17741a,a17742a,a17743a,a17746a,a17750a,a17751a,a17752a,a17755a,a17759a,a17760a,a17761a,a17764a,a17768a,a17769a,a17770a,a17773a,a17777a,a17778a,a17779a,a17782a,a17786a,a17787a,a17788a,a17791a,a17795a,a17796a,a17797a,a17800a,a17804a,a17805a,a17806a,a17809a,a17813a,a17814a,a17815a,a17818a,a17822a,a17823a,a17824a,a17827a,a17831a,a17832a,a17833a,a17836a,a17840a,a17841a,a17842a,a17845a,a17849a,a17850a,a17851a,a17854a,a17858a,a17859a,a17860a,a17863a,a17867a,a17868a,a17869a,a17872a,a17876a,a17877a,a17878a,a17881a,a17885a,a17886a,a17887a,a17890a,a17894a,a17895a,a17896a,a17899a,a17903a,a17904a,a17905a,a17908a,a17912a,a17913a,a17914a,a17917a,a17921a,a17922a,a17923a,a17926a,a17930a,a17931a,a17932a,a17935a,a17939a,a17940a,a17941a,a17944a,a17948a,a17949a,a17950a,a17953a,a17957a,a17958a,a17959a,a17962a,a17966a,a17967a,a17968a,a17971a,a17975a,a17976a,a17977a,a17980a,a17984a,a17985a,a17986a,a17989a,a17993a,a17994a,a17995a,a17998a,a18002a,a18003a,a18004a,a18007a,a18011a,a18012a,a18013a,a18016a,a18020a,a18021a,a18022a,a18025a,a18029a,a18030a,a18031a,a18034a,a18038a,a18039a,a18040a,a18043a,a18047a,a18048a,a18049a,a18052a,a18056a,a18057a,a18058a,a18061a,a18065a,a18066a,a18067a,a18070a,a18074a,a18075a,a18076a,a18079a,a18083a,a18084a,a18085a,a18088a,a18092a,a18093a,a18094a,a18097a,a18101a,a18102a,a18103a,a18106a,a18110a,a18111a,a18112a,a18115a,a18119a,a18120a,a18121a,a18124a,a18128a,a18129a,a18130a,a18133a,a18137a,a18138a,a18139a,a18142a,a18146a,a18147a,a18148a,a18151a,a18155a,a18156a,a18157a,a18160a,a18164a,a18165a,a18166a,a18169a,a18173a,a18174a,a18175a,a18178a,a18182a,a18183a,a18184a,a18187a,a18191a,a18192a,a18193a,a18196a,a18200a,a18201a,a18202a,a18205a,a18209a,a18210a,a18211a,a18214a,a18218a,a18219a,a18220a,a18223a,a18227a,a18228a,a18229a,a18232a,a18236a,a18237a,a18238a,a18241a,a18245a,a18246a,a18247a,a18250a,a18254a,a18255a,a18256a,a18259a,a18263a,a18264a,a18265a,a18268a,a18272a,a18273a,a18274a,a18277a,a18281a,a18282a,a18283a,a18286a,a18290a,a18291a,a18292a,a18295a,a18299a,a18300a,a18301a,a18304a,a18308a,a18309a,a18310a,a18313a,a18317a,a18318a,a18319a,a18322a,a18326a,a18327a,a18328a,a18331a,a18335a,a18336a,a18337a,a18340a,a18344a,a18345a,a18346a,a18349a,a18353a,a18354a,a18355a,a18358a,a18362a,a18363a,a18364a,a18367a,a18371a,a18372a,a18373a,a18376a,a18380a,a18381a,a18382a,a18385a,a18389a,a18390a,a18391a,a18394a,a18398a,a18399a,a18400a,a18403a,a18407a,a18408a,a18409a,a18412a,a18416a,a18417a,a18418a,a18421a,a18425a,a18426a,a18427a,a18430a,a18434a,a18435a,a18436a,a18439a,a18443a,a18444a,a18445a,a18448a,a18452a,a18453a,a18454a,a18457a,a18461a,a18462a,a18463a,a18466a,a18470a,a18471a,a18472a,a18475a,a18479a,a18480a,a18481a,a18484a,a18488a,a18489a,a18490a,a18493a,a18497a,a18498a,a18499a,a18502a,a18506a,a18507a,a18508a,a18511a,a18515a,a18516a,a18517a,a18520a,a18524a,a18525a,a18526a,a18529a,a18533a,a18534a,a18535a,a18538a,a18542a,a18543a,a18544a,a18547a,a18551a,a18552a,a18553a,a18556a,a18560a,a18561a,a18562a,a18565a,a18569a,a18570a,a18571a,a18574a,a18578a,a18579a,a18580a,a18583a,a18587a,a18588a,a18589a,a18592a,a18596a,a18597a,a18598a,a18601a,a18605a,a18606a,a18607a,a18610a,a18614a,a18615a,a18616a,a18619a,a18623a,a18624a,a18625a,a18628a,a18632a,a18633a,a18634a,a18637a,a18641a,a18642a,a18643a,a18646a,a18650a,a18651a,a18652a,a18655a,a18659a,a18660a,a18661a,a18664a,a18668a,a18669a,a18670a,a18673a,a18677a,a18678a,a18679a,a18682a,a18686a,a18687a,a18688a,a18691a,a18695a,a18696a,a18697a,a18700a,a18704a,a18705a,a18706a,a18709a,a18713a,a18714a,a18715a,a18718a,a18722a,a18723a,a18724a,a18727a,a18731a,a18732a,a18733a,a18736a,a18740a,a18741a,a18742a,a18745a,a18749a,a18750a,a18751a,a18754a,a18758a,a18759a,a18760a,a18763a,a18767a,a18768a,a18769a,a18772a,a18776a,a18777a,a18778a,a18781a,a18785a,a18786a,a18787a,a18790a,a18794a,a18795a,a18796a,a18799a,a18803a,a18804a,a18805a,a18808a,a18812a,a18813a,a18814a,a18817a,a18821a,a18822a,a18823a,a18826a,a18830a,a18831a,a18832a,a18835a,a18839a,a18840a,a18841a,a18844a,a18848a,a18849a,a18850a,a18853a,a18857a,a18858a,a18859a,a18862a,a18866a,a18867a,a18868a,a18871a,a18875a,a18876a,a18877a,a18880a,a18884a,a18885a,a18886a,a18889a,a18893a,a18894a,a18895a,a18898a,a18902a,a18903a,a18904a,a18907a,a18911a,a18912a,a18913a,a18916a,a18920a,a18921a,a18922a,a18925a,a18929a,a18930a,a18931a,a18934a,a18938a,a18939a,a18940a,a18943a,a18947a,a18948a,a18949a,a18952a,a18956a,a18957a,a18958a,a18961a,a18965a,a18966a,a18967a,a18970a,a18974a,a18975a,a18976a,a18979a,a18983a,a18984a,a18985a,a18988a,a18992a,a18993a,a18994a,a18997a,a19001a,a19002a,a19003a,a19006a,a19010a,a19011a,a19012a,a19015a,a19019a,a19020a,a19021a,a19024a,a19028a,a19029a,a19030a,a19033a,a19037a,a19038a,a19039a,a19042a,a19046a,a19047a,a19048a,a19051a,a19055a,a19056a,a19057a,a19060a,a19064a,a19065a,a19066a,a19069a,a19073a,a19074a,a19075a,a19078a,a19082a,a19083a,a19084a,a19087a,a19091a,a19092a,a19093a,a19096a,a19100a,a19101a,a19102a,a19105a,a19109a,a19110a,a19111a,a19114a,a19118a,a19119a,a19120a,a19123a,a19127a,a19128a,a19129a,a19132a,a19136a,a19137a,a19138a,a19141a,a19145a,a19146a,a19147a,a19150a,a19154a,a19155a,a19156a,a19159a,a19163a,a19164a,a19165a,a19168a,a19172a,a19173a,a19174a,a19177a,a19181a,a19182a,a19183a,a19186a,a19190a,a19191a,a19192a,a19195a,a19199a,a19200a,a19201a,a19204a,a19208a,a19209a,a19210a,a19213a,a19217a,a19218a,a19219a,a19222a,a19226a,a19227a,a19228a,a19231a,a19235a,a19236a,a19237a,a19240a,a19244a,a19245a,a19246a,a19249a,a19253a,a19254a,a19255a,a19258a,a19262a,a19263a,a19264a,a19267a,a19271a,a19272a,a19273a,a19276a,a19280a,a19281a,a19282a,a19285a,a19289a,a19290a,a19291a,a19294a,a19298a,a19299a,a19300a,a19303a,a19307a,a19308a,a19309a,a19312a,a19316a,a19317a,a19318a,a19321a,a19325a,a19326a,a19327a,a19330a,a19334a,a19335a,a19336a,a19339a,a19343a,a19344a,a19345a,a19348a,a19352a,a19353a,a19354a,a19357a,a19361a,a19362a,a19363a,a19366a,a19370a,a19371a,a19372a,a19375a,a19379a,a19380a,a19381a,a19384a,a19388a,a19389a,a19390a,a19393a,a19397a,a19398a,a19399a,a19402a,a19406a,a19407a,a19408a,a19411a,a19415a,a19416a,a19417a,a19420a,a19424a,a19425a,a19426a,a19429a,a19433a,a19434a,a19435a,a19438a,a19442a,a19443a,a19444a,a19447a,a19451a,a19452a,a19453a,a19456a,a19460a,a19461a,a19462a,a19465a,a19469a,a19470a,a19471a,a19474a,a19478a,a19479a,a19480a,a19483a,a19487a,a19488a,a19489a,a19492a,a19496a,a19497a,a19498a,a19501a,a19505a,a19506a,a19507a,a19510a,a19514a,a19515a,a19516a,a19519a,a19523a,a19524a,a19525a,a19528a,a19532a,a19533a,a19534a,a19537a,a19541a,a19542a,a19543a,a19546a,a19550a,a19551a,a19552a,a19555a,a19559a,a19560a,a19561a,a19564a,a19568a,a19569a,a19570a,a19573a,a19577a,a19578a,a19579a,a19582a,a19586a,a19587a,a19588a,a19591a,a19595a,a19596a,a19597a,a19600a,a19604a,a19605a,a19606a,a19609a,a19613a,a19614a,a19615a,a19618a,a19622a,a19623a,a19624a,a19627a,a19631a,a19632a,a19633a,a19636a,a19640a,a19641a,a19642a,a19645a,a19649a,a19650a,a19651a,a19654a,a19658a,a19659a,a19660a,a19663a,a19667a,a19668a,a19669a,a19672a,a19676a,a19677a,a19678a,a19681a,a19685a,a19686a,a19687a,a19690a,a19694a,a19695a,a19696a,a19699a,a19703a,a19704a,a19705a,a19708a,a19712a,a19713a,a19714a,a19717a,a19721a,a19722a,a19723a,a19726a,a19730a,a19731a,a19732a,a19735a,a19739a,a19740a,a19741a,a19744a,a19748a,a19749a,a19750a,a19753a,a19757a,a19758a,a19759a,a19762a,a19766a,a19767a,a19768a,a19771a,a19775a,a19776a,a19777a,a19780a,a19784a,a19785a,a19786a,a19789a,a19793a,a19794a,a19795a,a19798a,a19802a,a19803a,a19804a,a19807a,a19811a,a19812a,a19813a,a19816a,a19820a,a19821a,a19822a,a19825a,a19829a,a19830a,a19831a,a19834a,a19838a,a19839a,a19840a,a19843a,a19847a,a19848a,a19849a,a19852a,a19856a,a19857a,a19858a,a19861a,a19865a,a19866a,a19867a,a19870a,a19874a,a19875a,a19876a,a19879a,a19883a,a19884a,a19885a,a19888a,a19892a,a19893a,a19894a,a19897a,a19901a,a19902a,a19903a,a19906a,a19910a,a19911a,a19912a,a19915a,a19919a,a19920a,a19921a,a19924a,a19928a,a19929a,a19930a,a19933a,a19937a,a19938a,a19939a,a19942a,a19946a,a19947a,a19948a,a19951a,a19955a,a19956a,a19957a,a19960a,a19964a,a19965a,a19966a,a19969a,a19973a,a19974a,a19975a,a19978a,a19982a,a19983a,a19984a,a19987a,a19991a,a19992a,a19993a,a19996a,a20000a,a20001a,a20002a,a20005a,a20009a,a20010a,a20011a,a20014a,a20018a,a20019a,a20020a,a20023a,a20027a,a20028a,a20029a,a20032a,a20036a,a20037a,a20038a,a20041a,a20045a,a20046a,a20047a,a20050a,a20054a,a20055a,a20056a,a20059a,a20063a,a20064a,a20065a,a20068a,a20072a,a20073a,a20074a,a20077a,a20081a,a20082a,a20083a,a20086a,a20090a,a20091a,a20092a,a20095a,a20099a,a20100a,a20101a,a20104a,a20108a,a20109a,a20110a,a20113a,a20117a,a20118a,a20119a,a20122a,a20126a,a20127a,a20128a,a20131a,a20135a,a20136a,a20137a,a20140a,a20144a,a20145a,a20146a,a20149a,a20153a,a20154a,a20155a,a20158a,a20162a,a20163a,a20164a,a20167a,a20171a,a20172a,a20173a,a20176a,a20180a,a20181a,a20182a,a20185a,a20189a,a20190a,a20191a,a20194a,a20198a,a20199a,a20200a,a20203a,a20207a,a20208a,a20209a,a20212a,a20216a,a20217a,a20218a,a20221a,a20225a,a20226a,a20227a,a20230a,a20234a,a20235a,a20236a,a20239a,a20243a,a20244a,a20245a,a20248a,a20252a,a20253a,a20254a,a20257a,a20261a,a20262a,a20263a,a20266a,a20270a,a20271a,a20272a,a20275a,a20279a,a20280a,a20281a,a20284a,a20288a,a20289a,a20290a,a20293a,a20297a,a20298a,a20299a,a20302a,a20306a,a20307a,a20308a,a20311a,a20315a,a20316a,a20317a,a20320a,a20324a,a20325a,a20326a,a20329a,a20333a,a20334a,a20335a,a20338a,a20342a,a20343a,a20344a,a20347a,a20351a,a20352a,a20353a,a20356a,a20360a,a20361a,a20362a,a20365a,a20369a,a20370a,a20371a,a20374a,a20378a,a20379a,a20380a,a20383a,a20387a,a20388a,a20389a,a20392a,a20396a,a20397a,a20398a,a20401a,a20405a,a20406a,a20407a,a20410a,a20414a,a20415a,a20416a,a20419a,a20423a,a20424a,a20425a,a20428a,a20432a,a20433a,a20434a,a20437a,a20441a,a20442a,a20443a,a20446a,a20450a,a20451a,a20452a,a20455a,a20459a,a20460a,a20461a,a20464a,a20468a,a20469a,a20470a,a20473a,a20477a,a20478a,a20479a,a20482a,a20486a,a20487a,a20488a,a20491a,a20495a,a20496a,a20497a,a20500a,a20504a,a20505a,a20506a,a20509a,a20513a,a20514a,a20515a,a20518a,a20522a,a20523a,a20524a,a20527a,a20531a,a20532a,a20533a,a20536a,a20540a,a20541a,a20542a,a20545a,a20549a,a20550a,a20551a,a20554a,a20558a,a20559a,a20560a,a20563a,a20567a,a20568a,a20569a,a20572a,a20576a,a20577a,a20578a,a20581a,a20585a,a20586a,a20587a,a20590a,a20594a,a20595a,a20596a,a20599a,a20603a,a20604a,a20605a,a20608a,a20612a,a20613a,a20614a,a20617a,a20621a,a20622a,a20623a,a20626a,a20630a,a20631a,a20632a,a20635a,a20639a,a20640a,a20641a,a20644a,a20648a,a20649a,a20650a,a20653a,a20657a,a20658a,a20659a,a20662a,a20666a,a20667a,a20668a,a20671a,a20675a,a20676a,a20677a,a20680a,a20684a,a20685a,a20686a,a20689a,a20693a,a20694a,a20695a,a20698a,a20702a,a20703a,a20704a,a20707a,a20711a,a20712a,a20713a,a20716a,a20720a,a20721a,a20722a,a20725a,a20729a,a20730a,a20731a,a20734a,a20738a,a20739a,a20740a,a20743a,a20747a,a20748a,a20749a,a20752a,a20756a,a20757a,a20758a,a20761a,a20765a,a20766a,a20767a,a20770a,a20774a,a20775a,a20776a,a20779a,a20783a,a20784a,a20785a,a20788a,a20792a,a20793a,a20794a,a20797a,a20801a,a20802a,a20803a,a20806a,a20810a,a20811a,a20812a,a20815a,a20819a,a20820a,a20821a,a20824a,a20828a,a20829a,a20830a,a20833a,a20837a,a20838a,a20839a,a20842a,a20846a,a20847a,a20848a,a20851a,a20855a,a20856a,a20857a,a20860a,a20864a,a20865a,a20866a,a20869a,a20873a,a20874a,a20875a,a20878a,a20882a,a20883a,a20884a,a20887a,a20891a,a20892a,a20893a,a20896a,a20900a,a20901a,a20902a,a20905a,a20909a,a20910a,a20911a,a20914a,a20918a,a20919a,a20920a,a20923a,a20927a,a20928a,a20929a,a20932a,a20936a,a20937a,a20938a,a20941a,a20945a,a20946a,a20947a,a20950a,a20954a,a20955a,a20956a,a20959a,a20963a,a20964a,a20965a,a20968a,a20972a,a20973a,a20974a,a20977a,a20981a,a20982a,a20983a,a20986a,a20990a,a20991a,a20992a,a20995a,a20999a,a21000a,a21001a,a21004a,a21008a,a21009a,a21010a,a21013a,a21017a,a21018a,a21019a,a21022a,a21026a,a21027a,a21028a,a21031a,a21035a,a21036a,a21037a,a21040a,a21044a,a21045a,a21046a,a21049a,a21053a,a21054a,a21055a,a21058a,a21062a,a21063a,a21064a,a21067a,a21071a,a21072a,a21073a,a21076a,a21080a,a21081a,a21082a,a21085a,a21089a,a21090a,a21091a,a21094a,a21098a,a21099a,a21100a,a21103a,a21107a,a21108a,a21109a,a21112a,a21116a,a21117a,a21118a,a21121a,a21125a,a21126a,a21127a,a21130a,a21134a,a21135a,a21136a,a21139a,a21143a,a21144a,a21145a,a21148a,a21152a,a21153a,a21154a,a21157a,a21161a,a21162a,a21163a,a21166a,a21170a,a21171a,a21172a,a21175a,a21179a,a21180a,a21181a,a21184a,a21188a,a21189a,a21190a,a21193a,a21197a,a21198a,a21199a,a21202a,a21206a,a21207a,a21208a,a21211a,a21215a,a21216a,a21217a,a21220a,a21224a,a21225a,a21226a,a21229a,a21233a,a21234a,a21235a,a21238a,a21242a,a21243a,a21244a,a21247a,a21251a,a21252a,a21253a,a21256a,a21260a,a21261a,a21262a,a21265a,a21269a,a21270a,a21271a,a21274a,a21278a,a21279a,a21280a,a21283a,a21287a,a21288a,a21289a,a21292a,a21296a,a21297a,a21298a,a21301a,a21305a,a21306a,a21307a,a21310a,a21314a,a21315a,a21316a,a21319a,a21323a,a21324a,a21325a,a21328a,a21332a,a21333a,a21334a,a21337a,a21341a,a21342a,a21343a,a21346a,a21350a,a21351a,a21352a,a21355a,a21359a,a21360a,a21361a,a21364a,a21368a,a21369a,a21370a,a21373a,a21377a,a21378a,a21379a,a21382a,a21386a,a21387a,a21388a,a21391a,a21395a,a21396a,a21397a,a21400a,a21404a,a21405a,a21406a,a21409a,a21413a,a21414a,a21415a,a21418a,a21422a,a21423a,a21424a,a21427a,a21431a,a21432a,a21433a,a21436a,a21440a,a21441a,a21442a,a21445a,a21449a,a21450a,a21451a,a21454a,a21458a,a21459a,a21460a,a21463a,a21467a,a21468a,a21469a,a21472a,a21476a,a21477a,a21478a,a21481a,a21485a,a21486a,a21487a,a21490a,a21494a,a21495a,a21496a,a21499a,a21503a,a21504a,a21505a,a21508a,a21512a,a21513a,a21514a,a21517a,a21521a,a21522a,a21523a,a21526a,a21530a,a21531a,a21532a,a21535a,a21539a,a21540a,a21541a,a21544a,a21548a,a21549a,a21550a,a21553a,a21557a,a21558a,a21559a,a21562a,a21566a,a21567a,a21568a,a21571a,a21575a,a21576a,a21577a,a21580a,a21584a,a21585a,a21586a,a21589a,a21593a,a21594a,a21595a,a21598a,a21602a,a21603a,a21604a,a21607a,a21611a,a21612a,a21613a,a21616a,a21620a,a21621a,a21622a,a21625a,a21629a,a21630a,a21631a,a21634a,a21638a,a21639a,a21640a,a21643a,a21647a,a21648a,a21649a,a21652a,a21656a,a21657a,a21658a,a21661a,a21665a,a21666a,a21667a,a21670a,a21674a,a21675a,a21676a,a21679a,a21683a,a21684a,a21685a,a21688a,a21692a,a21693a,a21694a,a21697a,a21701a,a21702a,a21703a,a21706a,a21710a,a21711a,a21712a,a21715a,a21719a,a21720a,a21721a,a21724a,a21728a,a21729a,a21730a,a21733a,a21737a,a21738a,a21739a,a21742a,a21746a,a21747a,a21748a,a21751a,a21755a,a21756a,a21757a,a21760a,a21764a,a21765a,a21766a,a21769a,a21773a,a21774a,a21775a,a21778a,a21782a,a21783a,a21784a,a21787a,a21791a,a21792a,a21793a,a21796a,a21800a,a21801a,a21802a,a21805a,a21809a,a21810a,a21811a,a21814a,a21818a,a21819a,a21820a,a21823a,a21827a,a21828a,a21829a,a21832a,a21836a,a21837a,a21838a,a21841a,a21845a,a21846a,a21847a,a21850a,a21854a,a21855a,a21856a,a21859a,a21863a,a21864a,a21865a,a21868a,a21872a,a21873a,a21874a,a21877a,a21881a,a21882a,a21883a,a21886a,a21890a,a21891a,a21892a,a21895a,a21899a,a21900a,a21901a,a21904a,a21908a,a21909a,a21910a,a21913a,a21917a,a21918a,a21919a,a21922a,a21926a,a21927a,a21928a,a21931a,a21935a,a21936a,a21937a,a21940a,a21944a,a21945a,a21946a,a21949a,a21953a,a21954a,a21955a,a21958a,a21962a,a21963a,a21964a,a21967a,a21971a,a21972a,a21973a,a21976a,a21980a,a21981a,a21982a,a21985a,a21989a,a21990a,a21991a,a21994a,a21998a,a21999a,a22000a,a22003a,a22007a,a22008a,a22009a,a22012a,a22016a,a22017a,a22018a,a22021a,a22025a,a22026a,a22027a,a22030a,a22034a,a22035a,a22036a,a22039a,a22043a,a22044a,a22045a,a22048a,a22052a,a22053a,a22054a,a22057a,a22061a,a22062a,a22063a,a22066a,a22070a,a22071a,a22072a,a22075a,a22079a,a22080a,a22081a,a22084a,a22088a,a22089a,a22090a,a22093a,a22097a,a22098a,a22099a,a22102a,a22106a,a22107a,a22108a,a22111a,a22115a,a22116a,a22117a,a22120a,a22124a,a22125a,a22126a,a22129a,a22133a,a22134a,a22135a,a22138a,a22142a,a22143a,a22144a,a22147a,a22151a,a22152a,a22153a,a22156a,a22160a,a22161a,a22162a,a22165a,a22169a,a22170a,a22171a,a22174a,a22178a,a22179a,a22180a,a22183a,a22187a,a22188a,a22189a,a22192a,a22196a,a22197a,a22198a,a22201a,a22205a,a22206a,a22207a,a22210a,a22214a,a22215a,a22216a,a22219a,a22223a,a22224a,a22225a,a22228a,a22232a,a22233a,a22234a,a22237a,a22241a,a22242a,a22243a,a22246a,a22250a,a22251a,a22252a,a22255a,a22259a,a22260a,a22261a,a22264a,a22268a,a22269a,a22270a,a22273a,a22277a,a22278a,a22279a,a22282a,a22286a,a22287a,a22288a,a22291a,a22295a,a22296a,a22297a,a22300a,a22304a,a22305a,a22306a,a22309a,a22313a,a22314a,a22315a,a22318a,a22322a,a22323a,a22324a,a22327a,a22331a,a22332a,a22333a,a22336a,a22340a,a22341a,a22342a,a22345a,a22349a,a22350a,a22351a,a22354a,a22358a,a22359a,a22360a,a22363a,a22367a,a22368a,a22369a,a22372a,a22376a,a22377a,a22378a,a22381a,a22385a,a22386a,a22387a,a22390a,a22394a,a22395a,a22396a,a22399a,a22403a,a22404a,a22405a,a22408a,a22412a,a22413a,a22414a,a22417a,a22421a,a22422a,a22423a,a22426a,a22430a,a22431a,a22432a,a22435a,a22439a,a22440a,a22441a,a22444a,a22448a,a22449a,a22450a,a22453a,a22457a,a22458a,a22459a,a22462a,a22466a,a22467a,a22468a,a22471a,a22475a,a22476a,a22477a,a22480a,a22484a,a22485a,a22486a,a22489a,a22493a,a22494a,a22495a,a22498a,a22502a,a22503a,a22504a,a22507a,a22511a,a22512a,a22513a,a22516a,a22520a,a22521a,a22522a,a22525a,a22529a,a22530a,a22531a,a22534a,a22538a,a22539a,a22540a,a22543a,a22547a,a22548a,a22549a,a22552a,a22556a,a22557a,a22558a,a22561a,a22565a,a22566a,a22567a,a22570a,a22574a,a22575a,a22576a,a22579a,a22583a,a22584a,a22585a,a22588a,a22592a,a22593a,a22594a,a22597a,a22601a,a22602a,a22603a,a22606a,a22610a,a22611a,a22612a,a22615a,a22619a,a22620a,a22621a,a22624a,a22628a,a22629a,a22630a,a22633a,a22637a,a22638a,a22639a,a22642a,a22646a,a22647a,a22648a,a22651a,a22655a,a22656a,a22657a,a22660a,a22664a,a22665a,a22666a,a22669a,a22673a,a22674a,a22675a,a22678a,a22682a,a22683a,a22684a,a22687a,a22691a,a22692a,a22693a,a22696a,a22700a,a22701a,a22702a,a22705a,a22709a,a22710a,a22711a,a22714a,a22718a,a22719a,a22720a,a22723a,a22727a,a22728a,a22729a,a22733a,a22734a,a22738a,a22739a,a22740a,a22743a,a22747a,a22748a,a22749a,a22753a,a22754a,a22758a,a22759a,a22760a,a22763a,a22767a,a22768a,a22769a,a22773a,a22774a,a22778a,a22779a,a22780a,a22783a,a22787a,a22788a,a22789a,a22793a,a22794a,a22798a,a22799a,a22800a,a22803a,a22807a,a22808a,a22809a,a22813a,a22814a,a22818a,a22819a,a22820a,a22823a,a22827a,a22828a,a22829a,a22833a,a22834a,a22838a,a22839a,a22840a,a22843a,a22847a,a22848a,a22849a,a22853a,a22854a,a22858a,a22859a,a22860a,a22863a,a22867a,a22868a,a22869a,a22873a,a22874a,a22878a,a22879a,a22880a,a22883a,a22887a,a22888a,a22889a,a22893a,a22894a,a22898a,a22899a,a22900a,a22903a,a22907a,a22908a,a22909a,a22913a,a22914a,a22918a,a22919a,a22920a,a22923a,a22927a,a22928a,a22929a,a22933a,a22934a,a22938a,a22939a,a22940a,a22943a,a22947a,a22948a,a22949a,a22953a,a22954a,a22958a,a22959a,a22960a,a22963a,a22967a,a22968a,a22969a,a22973a,a22974a,a22978a,a22979a,a22980a,a22983a,a22987a,a22988a,a22989a,a22993a,a22994a,a22998a,a22999a,a23000a,a23003a,a23007a,a23008a,a23009a,a23013a,a23014a,a23018a,a23019a,a23020a,a23023a,a23027a,a23028a,a23029a,a23033a,a23034a,a23038a,a23039a,a23040a,a23043a,a23047a,a23048a,a23049a,a23053a,a23054a,a23058a,a23059a,a23060a,a23063a,a23067a,a23068a,a23069a,a23073a,a23074a,a23078a,a23079a,a23080a,a23083a,a23087a,a23088a,a23089a,a23093a,a23094a,a23098a,a23099a,a23100a,a23103a,a23107a,a23108a,a23109a,a23113a,a23114a,a23118a,a23119a,a23120a,a23123a,a23127a,a23128a,a23129a,a23133a,a23134a,a23138a,a23139a,a23140a,a23143a,a23147a,a23148a,a23149a,a23153a,a23154a,a23158a,a23159a,a23160a,a23163a,a23167a,a23168a,a23169a,a23173a,a23174a,a23178a,a23179a,a23180a,a23183a,a23187a,a23188a,a23189a,a23193a,a23194a,a23198a,a23199a,a23200a,a23203a,a23207a,a23208a,a23209a,a23213a,a23214a,a23218a,a23219a,a23220a,a23223a,a23227a,a23228a,a23229a,a23233a,a23234a,a23238a,a23239a,a23240a,a23243a,a23247a,a23248a,a23249a,a23253a,a23254a,a23258a,a23259a,a23260a,a23263a,a23267a,a23268a,a23269a,a23273a,a23274a,a23278a,a23279a,a23280a,a23283a,a23287a,a23288a,a23289a,a23293a,a23294a,a23298a,a23299a,a23300a,a23303a,a23307a,a23308a,a23309a,a23313a,a23314a,a23318a,a23319a,a23320a,a23323a,a23327a,a23328a,a23329a,a23333a,a23334a,a23338a,a23339a,a23340a,a23343a,a23347a,a23348a,a23349a,a23353a,a23354a,a23358a,a23359a,a23360a,a23363a,a23367a,a23368a,a23369a,a23373a,a23374a,a23378a,a23379a,a23380a,a23383a,a23387a,a23388a,a23389a,a23393a,a23394a,a23398a,a23399a,a23400a,a23403a,a23407a,a23408a,a23409a,a23413a,a23414a,a23418a,a23419a,a23420a,a23423a,a23427a,a23428a,a23429a,a23433a,a23434a,a23438a,a23439a,a23440a,a23443a,a23447a,a23448a,a23449a,a23453a,a23454a,a23458a,a23459a,a23460a,a23463a,a23467a,a23468a,a23469a,a23473a,a23474a,a23478a,a23479a,a23480a,a23483a,a23487a,a23488a,a23489a,a23493a,a23494a,a23498a,a23499a,a23500a,a23503a,a23507a,a23508a,a23509a,a23513a,a23514a,a23518a,a23519a,a23520a,a23523a,a23527a,a23528a,a23529a,a23533a,a23534a,a23538a,a23539a,a23540a,a23543a,a23547a,a23548a,a23549a,a23553a,a23554a,a23558a,a23559a,a23560a,a23563a,a23567a,a23568a,a23569a,a23573a,a23574a,a23578a,a23579a,a23580a,a23583a,a23587a,a23588a,a23589a,a23593a,a23594a,a23598a,a23599a,a23600a,a23603a,a23607a,a23608a,a23609a,a23613a,a23614a,a23618a,a23619a,a23620a,a23623a,a23627a,a23628a,a23629a,a23633a,a23634a,a23638a,a23639a,a23640a,a23643a,a23647a,a23648a,a23649a,a23653a,a23654a,a23658a,a23659a,a23660a,a23663a,a23667a,a23668a,a23669a,a23673a,a23674a,a23678a,a23679a,a23680a,a23683a,a23687a,a23688a,a23689a,a23693a,a23694a,a23698a,a23699a,a23700a,a23703a,a23707a,a23708a,a23709a,a23713a,a23714a,a23718a,a23719a,a23720a,a23723a,a23727a,a23728a,a23729a,a23733a,a23734a,a23738a,a23739a,a23740a,a23743a,a23747a,a23748a,a23749a,a23753a,a23754a,a23758a,a23759a,a23760a,a23763a,a23767a,a23768a,a23769a,a23773a,a23774a,a23778a,a23779a,a23780a,a23783a,a23787a,a23788a,a23789a,a23793a,a23794a,a23798a,a23799a,a23800a,a23803a,a23807a,a23808a,a23809a,a23813a,a23814a,a23818a,a23819a,a23820a,a23823a,a23827a,a23828a,a23829a,a23833a,a23834a,a23838a,a23839a,a23840a,a23843a,a23847a,a23848a,a23849a,a23853a,a23854a,a23858a,a23859a,a23860a,a23863a,a23867a,a23868a,a23869a,a23873a,a23874a,a23878a,a23879a,a23880a,a23883a,a23887a,a23888a,a23889a,a23893a,a23894a,a23898a,a23899a,a23900a,a23903a,a23907a,a23908a,a23909a,a23913a,a23914a,a23918a,a23919a,a23920a,a23923a,a23927a,a23928a,a23929a,a23933a,a23934a,a23938a,a23939a,a23940a,a23943a,a23947a,a23948a,a23949a,a23953a,a23954a,a23958a,a23959a,a23960a,a23963a,a23967a,a23968a,a23969a,a23973a,a23974a,a23978a,a23979a,a23980a,a23983a,a23987a,a23988a,a23989a,a23993a,a23994a,a23998a,a23999a,a24000a,a24003a,a24007a,a24008a,a24009a,a24013a,a24014a,a24018a,a24019a,a24020a,a24023a,a24027a,a24028a,a24029a,a24033a,a24034a,a24038a,a24039a,a24040a,a24043a,a24047a,a24048a,a24049a,a24053a,a24054a,a24058a,a24059a,a24060a,a24063a,a24067a,a24068a,a24069a,a24073a,a24074a,a24078a,a24079a,a24080a,a24083a,a24087a,a24088a,a24089a,a24093a,a24094a,a24098a,a24099a,a24100a,a24103a,a24107a,a24108a,a24109a,a24113a,a24114a,a24118a,a24119a,a24120a,a24123a,a24127a,a24128a,a24129a,a24133a,a24134a,a24138a,a24139a,a24140a,a24143a,a24147a,a24148a,a24149a,a24153a,a24154a,a24158a,a24159a,a24160a,a24163a,a24167a,a24168a,a24169a,a24173a,a24174a,a24178a,a24179a,a24180a,a24183a,a24187a,a24188a,a24189a,a24193a,a24194a,a24198a,a24199a,a24200a,a24203a,a24207a,a24208a,a24209a,a24213a,a24214a,a24218a,a24219a,a24220a,a24223a,a24227a,a24228a,a24229a,a24233a,a24234a,a24238a,a24239a,a24240a,a24243a,a24247a,a24248a,a24249a,a24253a,a24254a,a24258a,a24259a,a24260a,a24263a,a24267a,a24268a,a24269a,a24273a,a24274a,a24278a,a24279a,a24280a,a24283a,a24287a,a24288a,a24289a,a24293a,a24294a,a24298a,a24299a,a24300a,a24303a,a24307a,a24308a,a24309a,a24313a,a24314a,a24318a,a24319a,a24320a,a24323a,a24327a,a24328a,a24329a,a24333a,a24334a,a24338a,a24339a,a24340a,a24343a,a24347a,a24348a,a24349a,a24353a,a24354a,a24358a,a24359a,a24360a,a24363a,a24367a,a24368a,a24369a,a24373a,a24374a,a24378a,a24379a,a24380a,a24383a,a24387a,a24388a,a24389a,a24393a,a24394a,a24398a,a24399a,a24400a,a24403a,a24407a,a24408a,a24409a,a24413a,a24414a,a24418a,a24419a,a24420a,a24423a,a24427a,a24428a,a24429a,a24433a,a24434a,a24438a,a24439a,a24440a,a24443a,a24447a,a24448a,a24449a,a24453a,a24454a,a24458a,a24459a,a24460a,a24463a,a24467a,a24468a,a24469a,a24473a,a24474a,a24478a,a24479a,a24480a,a24483a,a24487a,a24488a,a24489a,a24493a,a24494a,a24498a,a24499a,a24500a,a24503a,a24507a,a24508a,a24509a,a24513a,a24514a,a24518a,a24519a,a24520a,a24523a,a24527a,a24528a,a24529a,a24533a,a24534a,a24538a,a24539a,a24540a,a24543a,a24547a,a24548a,a24549a,a24553a,a24554a,a24558a,a24559a,a24560a,a24563a,a24567a,a24568a,a24569a,a24573a,a24574a,a24578a,a24579a,a24580a,a24583a,a24587a,a24588a,a24589a,a24593a,a24594a,a24598a,a24599a,a24600a,a24603a,a24607a,a24608a,a24609a,a24613a,a24614a,a24618a,a24619a,a24620a,a24623a,a24627a,a24628a,a24629a,a24633a,a24634a,a24638a,a24639a,a24640a,a24643a,a24647a,a24648a,a24649a,a24653a,a24654a,a24658a,a24659a,a24660a,a24663a,a24667a,a24668a,a24669a,a24673a,a24674a,a24678a,a24679a,a24680a,a24683a,a24687a,a24688a,a24689a,a24693a,a24694a,a24698a,a24699a,a24700a,a24703a,a24707a,a24708a,a24709a,a24713a,a24714a,a24718a,a24719a,a24720a,a24723a,a24727a,a24728a,a24729a,a24733a,a24734a,a24738a,a24739a,a24740a,a24743a,a24747a,a24748a,a24749a,a24753a,a24754a,a24758a,a24759a,a24760a,a24763a,a24767a,a24768a,a24769a,a24773a,a24774a,a24778a,a24779a,a24780a,a24783a,a24787a,a24788a,a24789a,a24793a,a24794a,a24798a,a24799a,a24800a,a24803a,a24807a,a24808a,a24809a,a24813a,a24814a,a24818a,a24819a,a24820a,a24823a,a24827a,a24828a,a24829a,a24833a,a24834a,a24838a,a24839a,a24840a,a24843a,a24847a,a24848a,a24849a,a24853a,a24854a,a24858a,a24859a,a24860a,a24863a,a24867a,a24868a,a24869a,a24873a,a24874a,a24878a,a24879a,a24880a,a24883a,a24887a,a24888a,a24889a,a24893a,a24894a,a24898a,a24899a,a24900a,a24903a,a24907a,a24908a,a24909a,a24913a,a24914a,a24918a,a24919a,a24920a,a24923a,a24927a,a24928a,a24929a,a24933a,a24934a,a24938a,a24939a,a24940a,a24943a,a24947a,a24948a,a24949a,a24953a,a24954a,a24958a,a24959a,a24960a,a24963a,a24967a,a24968a,a24969a,a24973a,a24974a,a24978a,a24979a,a24980a,a24983a,a24987a,a24988a,a24989a,a24993a,a24994a,a24998a,a24999a,a25000a,a25003a,a25007a,a25008a,a25009a,a25013a,a25014a,a25018a,a25019a,a25020a,a25023a,a25027a,a25028a,a25029a,a25033a,a25034a,a25038a,a25039a,a25040a,a25043a,a25047a,a25048a,a25049a,a25053a,a25054a,a25058a,a25059a,a25060a,a25063a,a25067a,a25068a,a25069a,a25073a,a25074a,a25078a,a25079a,a25080a,a25083a,a25087a,a25088a,a25089a,a25093a,a25094a,a25098a,a25099a,a25100a,a25103a,a25107a,a25108a,a25109a,a25113a,a25114a,a25118a,a25119a,a25120a,a25123a,a25127a,a25128a,a25129a,a25133a,a25134a,a25138a,a25139a,a25140a,a25143a,a25147a,a25148a,a25149a,a25153a,a25154a,a25158a,a25159a,a25160a,a25163a,a25167a,a25168a,a25169a,a25173a,a25174a,a25178a,a25179a,a25180a,a25183a,a25187a,a25188a,a25189a,a25193a,a25194a,a25198a,a25199a,a25200a,a25203a,a25207a,a25208a,a25209a,a25213a,a25214a,a25218a,a25219a,a25220a,a25223a,a25227a,a25228a,a25229a,a25233a,a25234a,a25238a,a25239a,a25240a,a25243a,a25247a,a25248a,a25249a,a25253a,a25254a,a25258a,a25259a,a25260a,a25263a,a25267a,a25268a,a25269a,a25273a,a25274a,a25278a,a25279a,a25280a,a25283a,a25287a,a25288a,a25289a,a25293a,a25294a,a25298a,a25299a,a25300a,a25303a,a25307a,a25308a,a25309a,a25313a,a25314a,a25318a,a25319a,a25320a,a25323a,a25327a,a25328a,a25329a,a25333a,a25334a,a25338a,a25339a,a25340a,a25343a,a25347a,a25348a,a25349a,a25353a,a25354a,a25358a,a25359a,a25360a,a25363a,a25367a,a25368a,a25369a,a25373a,a25374a,a25378a,a25379a,a25380a,a25383a,a25387a,a25388a,a25389a,a25393a,a25394a,a25398a,a25399a,a25400a,a25403a,a25407a,a25408a,a25409a,a25413a,a25414a,a25418a,a25419a,a25420a,a25423a,a25427a,a25428a,a25429a,a25433a,a25434a,a25438a,a25439a,a25440a,a25443a,a25447a,a25448a,a25449a,a25453a,a25454a,a25458a,a25459a,a25460a,a25463a,a25467a,a25468a,a25469a,a25473a,a25474a,a25478a,a25479a,a25480a,a25483a,a25487a,a25488a,a25489a,a25493a,a25494a,a25498a,a25499a,a25500a,a25503a,a25507a,a25508a,a25509a,a25513a,a25514a,a25518a,a25519a,a25520a,a25523a,a25527a,a25528a,a25529a,a25533a,a25534a,a25538a,a25539a,a25540a,a25543a,a25547a,a25548a,a25549a,a25553a,a25554a,a25558a,a25559a,a25560a,a25563a,a25567a,a25568a,a25569a,a25573a,a25574a,a25578a,a25579a,a25580a,a25583a,a25587a,a25588a,a25589a,a25593a,a25594a,a25598a,a25599a,a25600a,a25603a,a25607a,a25608a,a25609a,a25613a,a25614a,a25618a,a25619a,a25620a,a25623a,a25627a,a25628a,a25629a,a25633a,a25634a,a25638a,a25639a,a25640a,a25643a,a25647a,a25648a,a25649a,a25653a,a25654a,a25658a,a25659a,a25660a,a25663a,a25667a,a25668a,a25669a,a25673a,a25674a,a25678a,a25679a,a25680a,a25683a,a25687a,a25688a,a25689a,a25693a,a25694a,a25698a,a25699a,a25700a,a25703a,a25707a,a25708a,a25709a,a25713a,a25714a,a25718a,a25719a,a25720a,a25723a,a25727a,a25728a,a25729a,a25733a,a25734a,a25738a,a25739a,a25740a,a25743a,a25747a,a25748a,a25749a,a25753a,a25754a,a25758a,a25759a,a25760a,a25763a,a25767a,a25768a,a25769a,a25773a,a25774a,a25778a,a25779a,a25780a,a25783a,a25787a,a25788a,a25789a,a25793a,a25794a,a25798a,a25799a,a25800a,a25803a,a25807a,a25808a,a25809a,a25813a,a25814a,a25818a,a25819a,a25820a,a25823a,a25827a,a25828a,a25829a,a25833a,a25834a,a25838a,a25839a,a25840a,a25843a,a25847a,a25848a,a25849a,a25853a,a25854a,a25858a,a25859a,a25860a,a25863a,a25867a,a25868a,a25869a,a25873a,a25874a,a25878a,a25879a,a25880a,a25883a,a25887a,a25888a,a25889a,a25893a,a25894a,a25898a,a25899a,a25900a,a25903a,a25907a,a25908a,a25909a,a25913a,a25914a,a25918a,a25919a,a25920a,a25923a,a25927a,a25928a,a25929a,a25933a,a25934a,a25938a,a25939a,a25940a,a25943a,a25947a,a25948a,a25949a,a25953a,a25954a,a25958a,a25959a,a25960a,a25963a,a25967a,a25968a,a25969a,a25973a,a25974a,a25978a,a25979a,a25980a,a25983a,a25987a,a25988a,a25989a,a25993a,a25994a,a25998a,a25999a,a26000a,a26003a,a26007a,a26008a,a26009a,a26013a,a26014a,a26018a,a26019a,a26020a,a26023a,a26027a,a26028a,a26029a,a26033a,a26034a,a26038a,a26039a,a26040a,a26043a,a26047a,a26048a,a26049a,a26053a,a26054a,a26058a,a26059a,a26060a,a26063a,a26067a,a26068a,a26069a,a26073a,a26074a,a26078a,a26079a,a26080a,a26083a,a26087a,a26088a,a26089a,a26093a,a26094a,a26098a,a26099a,a26100a,a26103a,a26107a,a26108a,a26109a,a26113a,a26114a,a26118a,a26119a,a26120a,a26123a,a26127a,a26128a,a26129a,a26133a,a26134a,a26138a,a26139a,a26140a,a26143a,a26147a,a26148a,a26149a,a26153a,a26154a,a26158a,a26159a,a26160a,a26163a,a26167a,a26168a,a26169a,a26173a,a26174a,a26178a,a26179a,a26180a,a26183a,a26187a,a26188a,a26189a,a26193a,a26194a,a26198a,a26199a,a26200a,a26203a,a26207a,a26208a,a26209a,a26213a,a26214a,a26218a,a26219a,a26220a,a26223a,a26227a,a26228a,a26229a,a26233a,a26234a,a26238a,a26239a,a26240a,a26243a,a26247a,a26248a,a26249a,a26253a,a26254a,a26258a,a26259a,a26260a,a26263a,a26267a,a26268a,a26269a,a26273a,a26274a,a26278a,a26279a,a26280a,a26283a,a26287a,a26288a,a26289a,a26293a,a26294a,a26298a,a26299a,a26300a,a26303a,a26307a,a26308a,a26309a,a26313a,a26314a,a26318a,a26319a,a26320a,a26323a,a26327a,a26328a,a26329a,a26333a,a26334a,a26338a,a26339a,a26340a,a26343a,a26347a,a26348a,a26349a,a26353a,a26354a,a26358a,a26359a,a26360a,a26363a,a26367a,a26368a,a26369a,a26373a,a26374a,a26378a,a26379a,a26380a,a26383a,a26387a,a26388a,a26389a,a26393a,a26394a,a26398a,a26399a,a26400a,a26403a,a26407a,a26408a,a26409a,a26413a,a26414a,a26418a,a26419a,a26420a,a26423a,a26427a,a26428a,a26429a,a26433a,a26434a,a26438a,a26439a,a26440a,a26443a,a26447a,a26448a,a26449a,a26453a,a26454a,a26458a,a26459a,a26460a,a26463a,a26467a,a26468a,a26469a,a26473a,a26474a,a26478a,a26479a,a26480a,a26483a,a26487a,a26488a,a26489a,a26493a,a26494a,a26498a,a26499a,a26500a,a26503a,a26507a,a26508a,a26509a,a26513a,a26514a,a26518a,a26519a,a26520a,a26523a,a26527a,a26528a,a26529a,a26533a,a26534a,a26538a,a26539a,a26540a,a26543a,a26547a,a26548a,a26549a,a26553a,a26554a,a26558a,a26559a,a26560a,a26563a,a26567a,a26568a,a26569a,a26573a,a26574a,a26578a,a26579a,a26580a,a26583a,a26587a,a26588a,a26589a,a26593a,a26594a,a26598a,a26599a,a26600a,a26603a,a26607a,a26608a,a26609a,a26613a,a26614a,a26618a,a26619a,a26620a,a26623a,a26627a,a26628a,a26629a,a26633a,a26634a,a26638a,a26639a,a26640a,a26643a,a26647a,a26648a,a26649a,a26653a,a26654a,a26658a,a26659a,a26660a,a26663a,a26667a,a26668a,a26669a,a26673a,a26674a,a26678a,a26679a,a26680a,a26683a,a26687a,a26688a,a26689a,a26693a,a26694a,a26698a,a26699a,a26700a,a26703a,a26707a,a26708a,a26709a,a26713a,a26714a,a26718a,a26719a,a26720a,a26723a,a26727a,a26728a,a26729a,a26733a,a26734a,a26738a,a26739a,a26740a,a26743a,a26747a,a26748a,a26749a,a26753a,a26754a,a26758a,a26759a,a26760a,a26763a,a26767a,a26768a,a26769a,a26773a,a26774a,a26778a,a26779a,a26780a,a26783a,a26787a,a26788a,a26789a,a26793a,a26794a,a26798a,a26799a,a26800a,a26803a,a26807a,a26808a,a26809a,a26813a,a26814a,a26818a,a26819a,a26820a,a26823a,a26827a,a26828a,a26829a,a26833a,a26834a,a26838a,a26839a,a26840a,a26843a,a26847a,a26848a,a26849a,a26853a,a26854a,a26858a,a26859a,a26860a,a26863a,a26867a,a26868a,a26869a,a26873a,a26874a,a26878a,a26879a,a26880a,a26883a,a26887a,a26888a,a26889a,a26893a,a26894a,a26898a,a26899a,a26900a,a26903a,a26907a,a26908a,a26909a,a26913a,a26914a,a26918a,a26919a,a26920a,a26923a,a26927a,a26928a,a26929a,a26933a,a26934a,a26938a,a26939a,a26940a,a26943a,a26947a,a26948a,a26949a,a26953a,a26954a,a26958a,a26959a,a26960a,a26963a,a26967a,a26968a,a26969a,a26973a,a26974a,a26978a,a26979a,a26980a,a26983a,a26987a,a26988a,a26989a,a26993a,a26994a,a26998a,a26999a,a27000a,a27003a,a27007a,a27008a,a27009a,a27013a,a27014a,a27018a,a27019a,a27020a,a27023a,a27027a,a27028a,a27029a,a27033a,a27034a,a27038a,a27039a,a27040a,a27043a,a27047a,a27048a,a27049a,a27053a,a27054a,a27058a,a27059a,a27060a,a27063a,a27067a,a27068a,a27069a,a27073a,a27074a,a27078a,a27079a,a27080a,a27083a,a27087a,a27088a,a27089a,a27093a,a27094a,a27098a,a27099a,a27100a,a27103a,a27107a,a27108a,a27109a,a27113a,a27114a,a27118a,a27119a,a27120a,a27123a,a27127a,a27128a,a27129a,a27133a,a27134a,a27138a,a27139a,a27140a,a27143a,a27147a,a27148a,a27149a,a27153a,a27154a,a27158a,a27159a,a27160a,a27163a,a27167a,a27168a,a27169a,a27173a,a27174a,a27178a,a27179a,a27180a,a27183a,a27187a,a27188a,a27189a,a27193a,a27194a,a27198a,a27199a,a27200a,a27203a,a27207a,a27208a,a27209a,a27213a,a27214a,a27218a,a27219a,a27220a,a27223a,a27227a,a27228a,a27229a,a27233a,a27234a,a27238a,a27239a,a27240a,a27243a,a27247a,a27248a,a27249a,a27253a,a27254a,a27258a,a27259a,a27260a,a27263a,a27267a,a27268a,a27269a,a27273a,a27274a,a27278a,a27279a,a27280a,a27283a,a27287a,a27288a,a27289a,a27293a,a27294a,a27298a,a27299a,a27300a,a27303a,a27307a,a27308a,a27309a,a27313a,a27314a,a27318a,a27319a,a27320a,a27323a,a27327a,a27328a,a27329a,a27333a,a27334a,a27338a,a27339a,a27340a,a27343a,a27347a,a27348a,a27349a,a27353a,a27354a,a27358a,a27359a,a27360a,a27363a,a27367a,a27368a,a27369a,a27373a,a27374a,a27378a,a27379a,a27380a,a27383a,a27387a,a27388a,a27389a,a27393a,a27394a,a27398a,a27399a,a27400a,a27403a,a27407a,a27408a,a27409a,a27413a,a27414a,a27418a,a27419a,a27420a,a27423a,a27427a,a27428a,a27429a,a27433a,a27434a,a27438a,a27439a,a27440a,a27443a,a27447a,a27448a,a27449a,a27453a,a27454a,a27458a,a27459a,a27460a,a27463a,a27467a,a27468a,a27469a,a27473a,a27474a,a27478a,a27479a,a27480a,a27483a,a27487a,a27488a,a27489a,a27493a,a27494a,a27498a,a27499a,a27500a,a27503a,a27507a,a27508a,a27509a,a27513a,a27514a,a27518a,a27519a,a27520a,a27523a,a27527a,a27528a,a27529a,a27533a,a27534a,a27538a,a27539a,a27540a,a27543a,a27547a,a27548a,a27549a,a27553a,a27554a,a27558a,a27559a,a27560a,a27563a,a27567a,a27568a,a27569a,a27573a,a27574a,a27578a,a27579a,a27580a,a27583a,a27587a,a27588a,a27589a,a27593a,a27594a,a27598a,a27599a,a27600a,a27603a,a27607a,a27608a,a27609a,a27613a,a27614a,a27618a,a27619a,a27620a,a27623a,a27627a,a27628a,a27629a,a27633a,a27634a,a27638a,a27639a,a27640a,a27643a,a27647a,a27648a,a27649a,a27653a,a27654a,a27658a,a27659a,a27660a,a27663a,a27667a,a27668a,a27669a,a27673a,a27674a,a27678a,a27679a,a27680a,a27683a,a27687a,a27688a,a27689a,a27693a,a27694a,a27698a,a27699a,a27700a,a27703a,a27707a,a27708a,a27709a,a27713a,a27714a,a27718a,a27719a,a27720a,a27723a,a27727a,a27728a,a27729a,a27733a,a27734a,a27738a,a27739a,a27740a,a27743a,a27747a,a27748a,a27749a,a27753a,a27754a,a27758a,a27759a,a27760a,a27763a,a27767a,a27768a,a27769a,a27773a,a27774a,a27778a,a27779a,a27780a,a27783a,a27787a,a27788a,a27789a,a27793a,a27794a,a27798a,a27799a,a27800a,a27803a,a27807a,a27808a,a27809a,a27813a,a27814a,a27818a,a27819a,a27820a,a27823a,a27827a,a27828a,a27829a,a27833a,a27834a,a27838a,a27839a,a27840a,a27843a,a27847a,a27848a,a27849a,a27853a,a27854a,a27858a,a27859a,a27860a,a27863a,a27867a,a27868a,a27869a,a27873a,a27874a,a27878a,a27879a,a27880a,a27883a,a27887a,a27888a,a27889a,a27893a,a27894a,a27898a,a27899a,a27900a,a27903a,a27907a,a27908a,a27909a,a27913a,a27914a,a27918a,a27919a,a27920a,a27923a,a27927a,a27928a,a27929a,a27933a,a27934a,a27938a,a27939a,a27940a,a27943a,a27947a,a27948a,a27949a,a27953a,a27954a,a27958a,a27959a,a27960a,a27963a,a27967a,a27968a,a27969a,a27973a,a27974a,a27978a,a27979a,a27980a,a27983a,a27987a,a27988a,a27989a,a27993a,a27994a,a27998a,a27999a,a28000a,a28003a,a28007a,a28008a,a28009a,a28013a,a28014a,a28018a,a28019a,a28020a,a28023a,a28027a,a28028a,a28029a,a28033a,a28034a,a28038a,a28039a,a28040a,a28043a,a28047a,a28048a,a28049a,a28053a,a28054a,a28058a,a28059a,a28060a,a28063a,a28067a,a28068a,a28069a,a28073a,a28074a,a28078a,a28079a,a28080a,a28083a,a28087a,a28088a,a28089a,a28093a,a28094a,a28098a,a28099a,a28100a,a28103a,a28107a,a28108a,a28109a,a28113a,a28114a,a28118a,a28119a,a28120a,a28123a,a28127a,a28128a,a28129a,a28133a,a28134a,a28138a,a28139a,a28140a,a28143a,a28147a,a28148a,a28149a,a28153a,a28154a,a28158a,a28159a,a28160a,a28163a,a28167a,a28168a,a28169a,a28173a,a28174a,a28178a,a28179a,a28180a,a28183a,a28187a,a28188a,a28189a,a28193a,a28194a,a28198a,a28199a,a28200a,a28203a,a28207a,a28208a,a28209a,a28213a,a28214a,a28218a,a28219a,a28220a,a28223a,a28227a,a28228a,a28229a,a28233a,a28234a,a28238a,a28239a,a28240a,a28243a,a28247a,a28248a,a28249a,a28253a,a28254a,a28258a,a28259a,a28260a,a28263a,a28267a,a28268a,a28269a,a28273a,a28274a,a28278a,a28279a,a28280a,a28283a,a28287a,a28288a,a28289a,a28293a,a28294a,a28298a,a28299a,a28300a,a28303a,a28307a,a28308a,a28309a,a28313a,a28314a,a28318a,a28319a,a28320a,a28323a,a28327a,a28328a,a28329a,a28333a,a28334a,a28338a,a28339a,a28340a,a28343a,a28347a,a28348a,a28349a,a28353a,a28354a,a28358a,a28359a,a28360a,a28363a,a28367a,a28368a,a28369a,a28373a,a28374a,a28378a,a28379a,a28380a,a28383a,a28387a,a28388a,a28389a,a28393a,a28394a,a28398a,a28399a,a28400a,a28403a,a28407a,a28408a,a28409a,a28413a,a28414a,a28418a,a28419a,a28420a,a28423a,a28427a,a28428a,a28429a,a28433a,a28434a,a28438a,a28439a,a28440a,a28443a,a28447a,a28448a,a28449a,a28453a,a28454a,a28458a,a28459a,a28460a,a28463a,a28467a,a28468a,a28469a,a28473a,a28474a,a28478a,a28479a,a28480a,a28483a,a28487a,a28488a,a28489a,a28493a,a28494a,a28498a,a28499a,a28500a,a28503a,a28507a,a28508a,a28509a,a28513a,a28514a,a28518a,a28519a,a28520a,a28523a,a28527a,a28528a,a28529a,a28533a,a28534a,a28538a,a28539a,a28540a,a28543a,a28547a,a28548a,a28549a,a28553a,a28554a,a28558a,a28559a,a28560a,a28563a,a28567a,a28568a,a28569a,a28573a,a28574a,a28578a,a28579a,a28580a,a28583a,a28587a,a28588a,a28589a,a28593a,a28594a,a28598a,a28599a,a28600a,a28603a,a28607a,a28608a,a28609a,a28613a,a28614a,a28618a,a28619a,a28620a,a28623a,a28627a,a28628a,a28629a,a28633a,a28634a,a28638a,a28639a,a28640a,a28643a,a28647a,a28648a,a28649a,a28653a,a28654a,a28658a,a28659a,a28660a,a28663a,a28667a,a28668a,a28669a,a28673a,a28674a,a28678a,a28679a,a28680a,a28683a,a28687a,a28688a,a28689a,a28693a,a28694a,a28698a,a28699a,a28700a,a28703a,a28707a,a28708a,a28709a,a28713a,a28714a,a28718a,a28719a,a28720a,a28723a,a28727a,a28728a,a28729a,a28733a,a28734a,a28738a,a28739a,a28740a,a28743a,a28747a,a28748a,a28749a,a28753a,a28754a,a28758a,a28759a,a28760a,a28763a,a28767a,a28768a,a28769a,a28773a,a28774a,a28778a,a28779a,a28780a,a28783a,a28787a,a28788a,a28789a,a28793a,a28794a,a28798a,a28799a,a28800a,a28803a,a28807a,a28808a,a28809a,a28813a,a28814a,a28818a,a28819a,a28820a,a28823a,a28827a,a28828a,a28829a,a28833a,a28834a,a28838a,a28839a,a28840a,a28843a,a28847a,a28848a,a28849a,a28853a,a28854a,a28858a,a28859a,a28860a,a28863a,a28867a,a28868a,a28869a,a28873a,a28874a,a28878a,a28879a,a28880a,a28883a,a28887a,a28888a,a28889a,a28893a,a28894a,a28898a,a28899a,a28900a,a28903a,a28907a,a28908a,a28909a,a28913a,a28914a,a28918a,a28919a,a28920a,a28923a,a28927a,a28928a,a28929a,a28933a,a28934a,a28938a,a28939a,a28940a,a28943a,a28947a,a28948a,a28949a,a28953a,a28954a,a28958a,a28959a,a28960a,a28963a,a28967a,a28968a,a28969a,a28973a,a28974a,a28978a,a28979a,a28980a,a28983a,a28987a,a28988a,a28989a,a28993a,a28994a,a28998a,a28999a,a29000a,a29003a,a29007a,a29008a,a29009a,a29013a,a29014a,a29018a,a29019a,a29020a,a29023a,a29027a,a29028a,a29029a,a29033a,a29034a,a29038a,a29039a,a29040a,a29043a,a29047a,a29048a,a29049a,a29053a,a29054a,a29058a,a29059a,a29060a,a29063a,a29067a,a29068a,a29069a,a29073a,a29074a,a29078a,a29079a,a29080a,a29083a,a29087a,a29088a,a29089a,a29093a,a29094a,a29098a,a29099a,a29100a,a29103a,a29107a,a29108a,a29109a,a29113a,a29114a,a29118a,a29119a,a29120a,a29123a,a29127a,a29128a,a29129a,a29133a,a29134a,a29138a,a29139a,a29140a,a29143a,a29147a,a29148a,a29149a,a29153a,a29154a,a29158a,a29159a,a29160a,a29163a,a29167a,a29168a,a29169a,a29173a,a29174a,a29178a,a29179a,a29180a,a29183a,a29187a,a29188a,a29189a,a29193a,a29194a,a29198a,a29199a,a29200a,a29203a,a29207a,a29208a,a29209a,a29213a,a29214a,a29218a,a29219a,a29220a,a29223a,a29227a,a29228a,a29229a,a29233a,a29234a,a29238a,a29239a,a29240a,a29243a,a29247a,a29248a,a29249a,a29253a,a29254a,a29258a,a29259a,a29260a,a29263a,a29267a,a29268a,a29269a,a29273a,a29274a,a29278a,a29279a,a29280a,a29283a,a29287a,a29288a,a29289a,a29293a,a29294a,a29298a,a29299a,a29300a,a29303a,a29307a,a29308a,a29309a,a29313a,a29314a,a29318a,a29319a,a29320a,a29323a,a29327a,a29328a,a29329a,a29333a,a29334a,a29338a,a29339a,a29340a,a29343a,a29347a,a29348a,a29349a,a29353a,a29354a,a29358a,a29359a,a29360a,a29363a,a29367a,a29368a,a29369a,a29373a,a29374a,a29378a,a29379a,a29380a,a29383a,a29387a,a29388a,a29389a,a29393a,a29394a,a29398a,a29399a,a29400a,a29403a,a29407a,a29408a,a29409a,a29413a,a29414a,a29418a,a29419a,a29420a,a29423a,a29427a,a29428a,a29429a,a29433a,a29434a,a29438a,a29439a,a29440a,a29444a,a29445a,a29449a,a29450a,a29451a,a29455a,a29456a,a29460a,a29461a,a29462a,a29466a,a29467a,a29471a,a29472a,a29473a,a29477a,a29478a,a29482a,a29483a,a29484a,a29488a,a29489a,a29493a,a29494a,a29495a,a29499a,a29500a,a29504a,a29505a,a29506a,a29510a,a29511a,a29515a,a29516a,a29517a,a29521a,a29522a,a29526a,a29527a,a29528a,a29532a,a29533a,a29537a,a29538a,a29539a,a29543a,a29544a,a29548a,a29549a,a29550a,a29554a,a29555a,a29559a,a29560a,a29561a,a29565a,a29566a,a29570a,a29571a,a29572a,a29576a,a29577a,a29581a,a29582a,a29583a,a29587a,a29588a,a29592a,a29593a,a29594a,a29598a,a29599a,a29603a,a29604a,a29605a,a29609a,a29610a,a29614a,a29615a,a29616a,a29620a,a29621a,a29625a,a29626a,a29627a,a29631a,a29632a,a29636a,a29637a,a29638a,a29642a,a29643a,a29647a,a29648a,a29649a,a29653a,a29654a,a29658a,a29659a,a29660a,a29664a,a29665a,a29669a,a29670a,a29671a,a29675a,a29676a,a29680a,a29681a,a29682a,a29686a,a29687a,a29691a,a29692a,a29693a,a29697a,a29698a,a29702a,a29703a,a29704a,a29708a,a29709a,a29713a,a29714a,a29715a,a29719a,a29720a,a29724a,a29725a,a29726a,a29730a,a29731a,a29735a,a29736a,a29737a,a29741a,a29742a,a29746a,a29747a,a29748a,a29752a,a29753a,a29757a,a29758a,a29759a,a29763a,a29764a,a29768a,a29769a,a29770a,a29774a,a29775a,a29779a,a29780a,a29781a,a29785a,a29786a,a29790a,a29791a,a29792a,a29796a,a29797a,a29801a,a29802a,a29803a,a29807a,a29808a,a29812a,a29813a,a29814a,a29818a,a29819a,a29823a,a29824a,a29825a,a29829a,a29830a,a29834a,a29835a,a29836a,a29840a,a29841a,a29845a,a29846a,a29847a,a29851a,a29852a,a29856a,a29857a,a29858a,a29862a,a29863a,a29867a,a29868a,a29869a,a29873a,a29874a,a29878a,a29879a,a29880a,a29884a,a29885a,a29889a,a29890a,a29891a,a29895a,a29896a,a29900a,a29901a,a29902a,a29906a,a29907a,a29911a,a29912a,a29913a,a29917a,a29918a,a29922a,a29923a,a29924a,a29928a,a29929a,a29933a,a29934a,a29935a,a29939a,a29940a,a29944a,a29945a,a29946a,a29950a,a29951a,a29955a,a29956a,a29957a,a29961a,a29962a,a29966a,a29967a,a29968a,a29972a,a29973a,a29977a,a29978a,a29979a,a29983a,a29984a,a29988a,a29989a,a29990a,a29994a,a29995a,a29999a,a30000a,a30001a,a30005a,a30006a,a30010a,a30011a,a30012a,a30016a,a30017a,a30021a,a30022a,a30023a,a30027a,a30028a,a30032a,a30033a,a30034a,a30038a,a30039a,a30043a,a30044a,a30045a,a30049a,a30050a,a30054a,a30055a,a30056a,a30060a,a30061a,a30065a,a30066a,a30067a,a30071a,a30072a,a30076a,a30077a,a30078a,a30082a,a30083a,a30087a,a30088a,a30089a,a30093a,a30094a,a30098a,a30099a,a30100a,a30104a,a30105a,a30109a,a30110a,a30111a,a30115a,a30116a,a30120a,a30121a,a30122a,a30126a,a30127a,a30131a,a30132a,a30133a,a30137a,a30138a,a30142a,a30143a,a30144a,a30148a,a30149a,a30153a,a30154a,a30155a,a30159a,a30160a,a30164a,a30165a,a30166a,a30170a,a30171a,a30175a,a30176a,a30177a,a30181a,a30182a,a30186a,a30187a,a30188a,a30192a,a30193a,a30197a,a30198a,a30199a,a30203a,a30204a,a30208a,a30209a,a30210a,a30214a,a30215a,a30219a,a30220a,a30221a,a30225a,a30226a,a30230a,a30231a,a30232a,a30236a,a30237a,a30241a,a30242a,a30243a,a30247a,a30248a,a30252a,a30253a,a30254a,a30258a,a30259a,a30263a,a30264a,a30265a,a30269a,a30270a,a30274a,a30275a,a30276a,a30280a,a30281a,a30285a,a30286a,a30287a,a30291a,a30292a,a30296a,a30297a,a30298a,a30302a,a30303a,a30307a,a30308a,a30309a,a30313a,a30314a,a30318a,a30319a,a30320a,a30324a,a30325a,a30329a,a30330a,a30331a,a30335a,a30336a,a30340a,a30341a,a30342a,a30346a,a30347a,a30351a,a30352a,a30353a,a30357a,a30358a,a30362a,a30363a,a30364a,a30368a,a30369a,a30373a,a30374a,a30375a,a30379a,a30380a,a30384a,a30385a,a30386a,a30390a,a30391a,a30395a,a30396a,a30397a,a30401a,a30402a,a30406a,a30407a,a30408a,a30412a,a30413a,a30417a,a30418a,a30419a,a30423a,a30424a,a30428a,a30429a,a30430a,a30434a,a30435a,a30439a,a30440a,a30441a,a30445a,a30446a,a30450a,a30451a,a30452a,a30456a,a30457a,a30461a,a30462a,a30463a,a30467a,a30468a,a30472a,a30473a,a30474a,a30478a,a30479a,a30483a,a30484a,a30485a,a30489a,a30490a,a30494a,a30495a,a30496a,a30500a,a30501a,a30505a,a30506a,a30507a,a30511a,a30512a,a30516a,a30517a,a30518a,a30522a,a30523a,a30527a,a30528a,a30529a,a30533a,a30534a,a30538a,a30539a,a30540a,a30544a,a30545a,a30549a,a30550a,a30551a,a30555a,a30556a,a30560a,a30561a,a30562a,a30566a,a30567a,a30571a,a30572a,a30573a,a30577a,a30578a,a30582a,a30583a,a30584a,a30588a,a30589a,a30593a,a30594a,a30595a,a30599a,a30600a,a30604a,a30605a,a30606a,a30610a,a30611a,a30615a,a30616a,a30617a,a30621a,a30622a,a30626a,a30627a,a30628a,a30632a,a30633a,a30637a,a30638a,a30639a,a30643a,a30644a,a30648a,a30649a,a30650a,a30654a,a30655a,a30659a,a30660a,a30661a,a30665a,a30666a,a30670a,a30671a,a30672a,a30676a,a30677a,a30681a,a30682a,a30683a,a30687a,a30688a,a30692a,a30693a,a30694a,a30698a,a30699a,a30703a,a30704a,a30705a,a30709a,a30710a,a30714a,a30715a,a30716a,a30720a,a30721a,a30725a,a30726a,a30727a,a30731a,a30732a,a30736a,a30737a,a30738a,a30742a,a30743a,a30747a,a30748a,a30749a,a30753a,a30754a,a30758a,a30759a,a30760a,a30764a,a30765a,a30769a,a30770a,a30771a,a30775a,a30776a,a30780a,a30781a,a30782a,a30786a,a30787a,a30791a,a30792a,a30793a,a30797a,a30798a,a30802a,a30803a,a30804a,a30808a,a30809a,a30813a,a30814a,a30815a,a30819a,a30820a,a30824a,a30825a,a30826a,a30830a,a30831a,a30835a,a30836a,a30837a,a30841a,a30842a,a30846a,a30847a,a30848a,a30852a,a30853a,a30857a,a30858a,a30859a,a30863a,a30864a,a30868a,a30869a,a30870a,a30874a,a30875a,a30879a,a30880a,a30881a,a30885a,a30886a,a30890a,a30891a,a30892a,a30896a,a30897a,a30901a,a30902a,a30903a,a30907a,a30908a,a30912a,a30913a,a30914a,a30918a,a30919a,a30923a,a30924a,a30925a,a30929a,a30930a,a30934a,a30935a,a30936a,a30940a,a30941a,a30945a,a30946a,a30947a,a30951a,a30952a,a30956a,a30957a,a30958a,a30962a,a30963a,a30967a,a30968a,a30969a,a30973a,a30974a,a30978a,a30979a,a30980a,a30984a,a30985a,a30989a,a30990a,a30991a,a30995a,a30996a,a31000a,a31001a,a31002a,a31006a,a31007a,a31011a,a31012a,a31013a,a31017a,a31018a,a31022a,a31023a,a31024a,a31028a,a31029a,a31033a,a31034a,a31035a,a31039a,a31040a,a31044a,a31045a,a31046a,a31050a,a31051a,a31055a,a31056a,a31057a,a31061a,a31062a,a31066a,a31067a,a31068a,a31072a,a31073a,a31077a,a31078a,a31079a,a31083a,a31084a,a31088a,a31089a,a31090a,a31094a,a31095a,a31099a,a31100a,a31101a,a31105a,a31106a,a31110a,a31111a,a31112a,a31116a,a31117a,a31121a,a31122a,a31123a,a31127a,a31128a,a31132a,a31133a,a31134a,a31138a,a31139a,a31143a,a31144a,a31145a,a31149a,a31150a,a31154a,a31155a,a31156a,a31160a,a31161a,a31165a,a31166a,a31167a,a31171a,a31172a,a31176a,a31177a,a31178a,a31182a,a31183a,a31187a,a31188a,a31189a,a31193a,a31194a,a31198a,a31199a,a31200a,a31204a,a31205a,a31209a,a31210a,a31211a,a31215a,a31216a,a31220a,a31221a,a31222a,a31226a,a31227a,a31231a,a31232a,a31233a,a31237a,a31238a,a31242a,a31243a,a31244a,a31248a,a31249a,a31253a,a31254a,a31255a,a31259a,a31260a,a31264a,a31265a,a31266a,a31270a,a31271a,a31275a,a31276a,a31277a,a31281a,a31282a,a31286a,a31287a,a31288a,a31292a,a31293a,a31297a,a31298a,a31299a,a31303a,a31304a,a31308a,a31309a,a31310a,a31314a,a31315a,a31319a,a31320a,a31321a,a31325a,a31326a,a31330a,a31331a,a31332a,a31336a,a31337a,a31341a,a31342a,a31343a,a31347a,a31348a,a31352a,a31353a,a31354a,a31358a,a31359a,a31363a,a31364a,a31365a,a31369a,a31370a,a31374a,a31375a,a31376a,a31380a,a31381a,a31385a,a31386a,a31387a,a31391a,a31392a,a31396a,a31397a,a31398a,a31402a,a31403a,a31407a,a31408a,a31409a,a31413a,a31414a,a31418a,a31419a,a31420a,a31424a,a31425a,a31429a,a31430a,a31431a,a31435a,a31436a,a31440a,a31441a,a31442a,a31446a,a31447a,a31451a,a31452a,a31453a,a31457a,a31458a,a31462a,a31463a,a31464a,a31468a,a31469a,a31473a,a31474a,a31475a,a31479a,a31480a,a31484a,a31485a,a31486a,a31490a,a31491a,a31495a,a31496a,a31497a,a31501a,a31502a,a31506a,a31507a,a31508a,a31512a,a31513a,a31517a,a31518a,a31519a,a31523a,a31524a,a31528a,a31529a,a31530a,a31534a,a31535a,a31539a,a31540a,a31541a,a31545a,a31546a,a31550a,a31551a,a31552a,a31556a,a31557a,a31561a,a31562a,a31563a,a31567a,a31568a,a31572a,a31573a,a31574a,a31578a,a31579a,a31583a,a31584a,a31585a,a31589a,a31590a,a31594a,a31595a,a31596a,a31600a,a31601a,a31605a,a31606a,a31607a,a31611a,a31612a,a31616a,a31617a,a31618a,a31622a,a31623a,a31627a,a31628a,a31629a,a31633a,a31634a,a31638a,a31639a,a31640a,a31644a,a31645a,a31649a,a31650a,a31651a,a31655a,a31656a,a31660a,a31661a,a31662a,a31666a,a31667a,a31671a,a31672a,a31673a,a31677a,a31678a,a31682a,a31683a,a31684a,a31688a,a31689a,a31693a,a31694a,a31695a,a31699a,a31700a,a31704a,a31705a,a31706a,a31710a,a31711a,a31715a,a31716a,a31717a,a31721a,a31722a,a31726a,a31727a,a31728a,a31732a,a31733a,a31737a,a31738a,a31739a,a31743a,a31744a,a31748a,a31749a,a31750a,a31754a,a31755a,a31759a,a31760a,a31761a,a31765a,a31766a,a31770a,a31771a,a31772a,a31776a,a31777a,a31781a,a31782a,a31783a,a31787a,a31788a,a31792a,a31793a,a31794a,a31798a,a31799a,a31803a,a31804a,a31805a,a31809a,a31810a,a31814a,a31815a,a31816a,a31820a,a31821a,a31825a,a31826a,a31827a,a31831a,a31832a,a31836a,a31837a,a31838a,a31842a,a31843a,a31847a,a31848a,a31849a,a31853a,a31854a,a31858a,a31859a,a31860a,a31864a,a31865a,a31869a,a31870a,a31871a,a31875a,a31876a,a31880a,a31881a,a31882a,a31886a,a31887a,a31891a,a31892a,a31893a,a31897a,a31898a,a31902a,a31903a,a31904a,a31908a,a31909a,a31913a,a31914a,a31915a,a31919a,a31920a,a31924a,a31925a,a31926a,a31930a,a31931a,a31935a,a31936a,a31937a,a31941a,a31942a,a31946a,a31947a,a31948a,a31952a,a31953a,a31957a,a31958a,a31959a,a31963a,a31964a,a31968a,a31969a,a31970a,a31974a,a31975a,a31979a,a31980a,a31981a,a31985a,a31986a,a31990a,a31991a,a31992a,a31996a,a31997a,a32001a,a32002a,a32003a,a32007a,a32008a,a32012a,a32013a,a32014a,a32018a,a32019a,a32023a,a32024a,a32025a,a32029a,a32030a,a32034a,a32035a,a32036a,a32040a,a32041a,a32045a,a32046a,a32047a,a32051a,a32052a,a32056a,a32057a,a32058a,a32062a,a32063a,a32067a,a32068a,a32069a,a32073a,a32074a,a32078a,a32079a,a32080a,a32084a,a32085a,a32089a,a32090a,a32091a,a32095a,a32096a,a32100a,a32101a,a32102a,a32106a,a32107a,a32111a,a32112a,a32113a,a32117a,a32118a,a32122a,a32123a,a32124a,a32128a,a32129a,a32133a,a32134a,a32135a,a32139a,a32140a,a32144a,a32145a,a32146a,a32150a,a32151a,a32155a,a32156a,a32157a,a32161a,a32162a,a32166a,a32167a,a32168a,a32172a,a32173a,a32177a,a32178a,a32179a,a32183a,a32184a,a32188a,a32189a,a32190a,a32194a,a32195a,a32199a,a32200a,a32201a,a32205a,a32206a,a32210a,a32211a,a32212a,a32216a,a32217a,a32221a,a32222a,a32223a,a32227a,a32228a,a32232a,a32233a,a32234a,a32238a,a32239a,a32243a,a32244a,a32245a,a32249a,a32250a,a32254a,a32255a,a32256a,a32260a,a32261a,a32265a,a32266a,a32267a,a32271a,a32272a,a32276a,a32277a,a32278a,a32282a,a32283a,a32287a,a32288a,a32289a,a32293a,a32294a,a32298a,a32299a,a32300a,a32304a,a32305a,a32309a,a32310a,a32311a,a32315a,a32316a,a32320a,a32321a,a32322a,a32326a,a32327a,a32331a,a32332a,a32333a,a32337a,a32338a,a32342a,a32343a,a32344a,a32348a,a32349a,a32353a,a32354a,a32355a,a32359a,a32360a,a32364a,a32365a,a32366a,a32370a,a32371a,a32375a,a32376a,a32377a,a32381a,a32382a,a32386a,a32387a,a32388a,a32392a,a32393a,a32397a,a32398a,a32399a,a32403a,a32404a,a32408a,a32409a,a32410a,a32414a,a32415a,a32419a,a32420a,a32421a,a32425a,a32426a,a32430a,a32431a,a32432a,a32436a,a32437a,a32441a,a32442a,a32443a,a32447a,a32448a,a32452a,a32453a,a32454a,a32458a,a32459a,a32463a,a32464a,a32465a,a32469a,a32470a,a32474a,a32475a,a32476a,a32480a,a32481a,a32485a,a32486a,a32487a,a32491a,a32492a,a32496a,a32497a,a32498a,a32502a,a32503a,a32507a,a32508a,a32509a,a32513a,a32514a,a32518a,a32519a,a32520a,a32524a,a32525a,a32529a,a32530a,a32531a,a32535a,a32536a,a32540a,a32541a,a32542a,a32546a,a32547a,a32551a,a32552a,a32553a,a32557a,a32558a,a32562a,a32563a,a32564a,a32568a,a32569a,a32573a,a32574a,a32575a,a32579a,a32580a,a32584a,a32585a,a32586a,a32590a,a32591a,a32595a,a32596a,a32597a,a32601a,a32602a,a32606a,a32607a,a32608a,a32612a,a32613a,a32617a,a32618a,a32619a,a32623a,a32624a,a32628a,a32629a,a32630a,a32634a,a32635a,a32639a,a32640a,a32641a,a32645a,a32646a,a32650a,a32651a,a32652a,a32656a,a32657a,a32661a,a32662a,a32663a,a32667a,a32668a,a32672a,a32673a,a32674a,a32678a,a32679a,a32683a,a32684a,a32685a,a32689a,a32690a,a32694a,a32695a,a32696a,a32700a,a32701a,a32705a,a32706a,a32707a,a32711a,a32712a,a32716a,a32717a,a32718a,a32722a,a32723a,a32727a,a32728a,a32729a,a32733a,a32734a,a32738a,a32739a,a32740a,a32744a,a32745a,a32749a,a32750a,a32751a,a32755a,a32756a,a32760a,a32761a,a32762a,a32766a,a32767a,a32771a,a32772a,a32773a,a32777a,a32778a,a32782a,a32783a,a32784a,a32788a,a32789a,a32793a,a32794a,a32795a,a32799a,a32800a,a32804a,a32805a,a32806a,a32810a,a32811a,a32815a,a32816a,a32817a,a32821a,a32822a,a32826a,a32827a,a32828a,a32832a,a32833a,a32837a,a32838a,a32839a,a32843a,a32844a,a32848a,a32849a,a32850a,a32854a,a32855a,a32859a,a32860a,a32861a,a32865a,a32866a,a32870a,a32871a,a32872a,a32876a,a32877a,a32881a,a32882a,a32883a,a32887a,a32888a,a32892a,a32893a,a32894a,a32898a,a32899a,a32903a,a32904a,a32905a,a32909a,a32910a,a32914a,a32915a,a32916a,a32920a,a32921a,a32925a,a32926a,a32927a,a32931a,a32932a,a32936a,a32937a,a32938a,a32942a,a32943a,a32947a,a32948a,a32949a,a32953a,a32954a,a32958a,a32959a,a32960a,a32964a,a32965a,a32969a,a32970a,a32971a,a32975a,a32976a,a32979a,a32982a,a32983a,a32984a,a32988a,a32989a,a32993a,a32994a,a32995a,a32999a,a33000a,a33003a,a33006a,a33007a,a33008a,a33012a,a33013a,a33017a,a33018a,a33019a,a33023a,a33024a,a33027a,a33030a,a33031a,a33032a,a33036a,a33037a,a33041a,a33042a,a33043a,a33047a,a33048a,a33051a,a33054a,a33055a,a33056a,a33060a,a33061a,a33065a,a33066a,a33067a,a33071a,a33072a,a33075a,a33078a,a33079a,a33080a,a33084a,a33085a,a33089a,a33090a,a33091a,a33095a,a33096a,a33099a,a33102a,a33103a,a33104a,a33108a,a33109a,a33113a,a33114a,a33115a,a33119a,a33120a,a33123a,a33126a,a33127a,a33128a,a33132a,a33133a,a33137a,a33138a,a33139a,a33143a,a33144a,a33147a,a33150a,a33151a,a33152a,a33156a,a33157a,a33161a,a33162a,a33163a,a33167a,a33168a,a33171a,a33174a,a33175a,a33176a,a33180a,a33181a,a33185a,a33186a,a33187a,a33191a,a33192a,a33195a,a33198a,a33199a,a33200a,a33204a,a33205a,a33209a,a33210a,a33211a,a33215a,a33216a,a33219a,a33222a,a33223a,a33224a,a33228a,a33229a,a33233a,a33234a,a33235a,a33239a,a33240a,a33243a,a33246a,a33247a,a33248a,a33252a,a33253a,a33257a,a33258a,a33259a,a33263a,a33264a,a33267a,a33270a,a33271a,a33272a,a33276a,a33277a,a33281a,a33282a,a33283a,a33287a,a33288a,a33291a,a33294a,a33295a,a33296a,a33300a,a33301a,a33305a,a33306a,a33307a,a33311a,a33312a,a33315a,a33318a,a33319a,a33320a,a33324a,a33325a,a33329a,a33330a,a33331a,a33335a,a33336a,a33339a,a33342a,a33343a,a33344a,a33348a,a33349a,a33353a,a33354a,a33355a,a33359a,a33360a,a33363a,a33366a,a33367a,a33368a,a33372a,a33373a,a33377a,a33378a,a33379a,a33383a,a33384a,a33387a,a33390a,a33391a,a33392a,a33396a,a33397a,a33401a,a33402a,a33403a,a33407a,a33408a,a33411a,a33414a,a33415a,a33416a,a33420a,a33421a,a33425a,a33426a,a33427a,a33431a,a33432a,a33435a,a33438a,a33439a,a33440a,a33444a,a33445a,a33449a,a33450a,a33451a,a33455a,a33456a,a33459a,a33462a,a33463a,a33464a,a33468a,a33469a,a33473a,a33474a,a33475a,a33479a,a33480a,a33483a,a33486a,a33487a,a33488a,a33492a,a33493a,a33497a,a33498a,a33499a,a33503a,a33504a,a33507a,a33510a,a33511a,a33512a,a33516a,a33517a,a33521a,a33522a,a33523a,a33527a,a33528a,a33531a,a33534a,a33535a,a33536a,a33540a,a33541a,a33545a,a33546a,a33547a,a33551a,a33552a,a33555a,a33558a,a33559a,a33560a,a33564a,a33565a,a33569a,a33570a,a33571a,a33575a,a33576a,a33579a,a33582a,a33583a,a33584a,a33588a,a33589a,a33593a,a33594a,a33595a,a33599a,a33600a,a33603a,a33606a,a33607a,a33608a,a33612a,a33613a,a33617a,a33618a,a33619a,a33623a,a33624a,a33627a,a33630a,a33631a,a33632a,a33636a,a33637a,a33641a,a33642a,a33643a,a33647a,a33648a,a33651a,a33654a,a33655a,a33656a,a33660a,a33661a,a33665a,a33666a,a33667a,a33671a,a33672a,a33675a,a33678a,a33679a,a33680a,a33684a,a33685a,a33689a,a33690a,a33691a,a33695a,a33696a,a33699a,a33702a,a33703a,a33704a,a33708a,a33709a,a33713a,a33714a,a33715a,a33719a,a33720a,a33723a,a33726a,a33727a,a33728a,a33732a,a33733a,a33737a,a33738a,a33739a,a33743a,a33744a,a33747a,a33750a,a33751a,a33752a,a33756a,a33757a,a33761a,a33762a,a33763a,a33767a,a33768a,a33771a,a33774a,a33775a,a33776a,a33780a,a33781a,a33785a,a33786a,a33787a,a33791a,a33792a,a33795a,a33798a,a33799a,a33800a,a33804a,a33805a,a33809a,a33810a,a33811a,a33815a,a33816a,a33819a,a33822a,a33823a,a33824a,a33828a,a33829a,a33833a,a33834a,a33835a,a33839a,a33840a,a33843a,a33846a,a33847a,a33848a,a33852a,a33853a,a33857a,a33858a,a33859a,a33863a,a33864a,a33867a,a33870a,a33871a,a33872a,a33876a,a33877a,a33881a,a33882a,a33883a,a33887a,a33888a,a33891a,a33894a,a33895a,a33896a,a33900a,a33901a,a33905a,a33906a,a33907a,a33911a,a33912a,a33915a,a33918a,a33919a,a33920a,a33924a,a33925a,a33929a,a33930a,a33931a,a33935a,a33936a,a33939a,a33942a,a33943a,a33944a,a33948a,a33949a,a33953a,a33954a,a33955a,a33959a,a33960a,a33963a,a33966a,a33967a,a33968a,a33972a,a33973a,a33977a,a33978a,a33979a,a33983a,a33984a,a33987a,a33990a,a33991a,a33992a,a33996a,a33997a,a34001a,a34002a,a34003a,a34007a,a34008a,a34011a,a34014a,a34015a,a34016a,a34020a,a34021a,a34025a,a34026a,a34027a,a34031a,a34032a,a34035a,a34038a,a34039a,a34040a,a34044a,a34045a,a34049a,a34050a,a34051a,a34055a,a34056a,a34059a,a34062a,a34063a,a34064a,a34068a,a34069a,a34073a,a34074a,a34075a,a34079a,a34080a,a34083a,a34086a,a34087a,a34088a,a34092a,a34093a,a34097a,a34098a,a34099a,a34103a,a34104a,a34107a,a34110a,a34111a,a34112a,a34116a,a34117a,a34121a,a34122a,a34123a,a34127a,a34128a,a34131a,a34134a,a34135a,a34136a,a34140a,a34141a,a34145a,a34146a,a34147a,a34151a,a34152a,a34155a,a34158a,a34159a,a34160a,a34164a,a34165a,a34169a,a34170a,a34171a,a34175a,a34176a,a34179a,a34182a,a34183a,a34184a,a34188a,a34189a,a34193a,a34194a,a34195a,a34199a,a34200a,a34203a,a34206a,a34207a,a34208a,a34212a,a34213a,a34217a,a34218a,a34219a,a34223a,a34224a,a34227a,a34230a,a34231a,a34232a,a34236a,a34237a,a34241a,a34242a,a34243a,a34247a,a34248a,a34251a,a34254a,a34255a,a34256a,a34260a,a34261a,a34265a,a34266a,a34267a,a34271a,a34272a,a34275a,a34278a,a34279a,a34280a,a34284a,a34285a,a34289a,a34290a,a34291a,a34295a,a34296a,a34299a,a34302a,a34303a,a34304a,a34308a,a34309a,a34313a,a34314a,a34315a,a34319a,a34320a,a34323a,a34326a,a34327a,a34328a,a34332a,a34333a,a34337a,a34338a,a34339a,a34343a,a34344a,a34347a,a34350a,a34351a,a34352a,a34356a,a34357a,a34361a,a34362a,a34363a,a34367a,a34368a,a34371a,a34374a,a34375a,a34376a,a34380a,a34381a,a34385a,a34386a,a34387a,a34391a,a34392a,a34395a,a34398a,a34399a,a34400a,a34404a,a34405a,a34409a,a34410a,a34411a,a34415a,a34416a,a34419a,a34422a,a34423a,a34424a,a34428a,a34429a,a34433a,a34434a,a34435a,a34439a,a34440a,a34443a,a34446a,a34447a,a34448a,a34452a,a34453a,a34457a,a34458a,a34459a,a34463a,a34464a,a34467a,a34470a,a34471a,a34472a,a34476a,a34477a,a34481a,a34482a,a34483a,a34487a,a34488a,a34491a,a34494a,a34495a,a34496a,a34500a,a34501a,a34504a,a34507a,a34508a,a34509a,a34513a,a34514a,a34517a,a34520a,a34521a,a34522a,a34526a,a34527a,a34530a,a34533a,a34534a,a34535a,a34539a,a34540a,a34543a,a34546a,a34547a,a34548a,a34552a,a34553a,a34556a,a34559a,a34560a,a34561a,a34565a,a34566a,a34569a,a34572a,a34573a,a34574a,a34578a,a34579a,a34582a,a34585a,a34586a,a34587a,a34591a,a34592a,a34595a,a34598a,a34599a,a34600a,a34604a,a34605a,a34608a,a34611a,a34612a,a34613a,a34617a,a34618a,a34621a,a34624a,a34625a,a34626a,a34630a,a34631a,a34634a,a34637a,a34638a,a34639a,a34643a,a34644a,a34647a,a34650a,a34651a,a34652a,a34656a,a34657a,a34660a,a34663a,a34664a,a34665a,a34669a,a34670a,a34673a,a34676a,a34677a,a34678a,a34682a,a34683a,a34686a,a34689a,a34690a,a34691a,a34695a,a34696a,a34699a,a34702a,a34703a,a34704a,a34708a,a34709a,a34712a,a34715a,a34716a,a34717a,a34721a,a34722a,a34725a,a34728a,a34729a,a34730a,a34734a,a34735a,a34738a,a34741a,a34742a,a34743a,a34747a,a34748a,a34751a,a34754a,a34755a,a34756a,a34760a,a34761a,a34764a,a34767a,a34768a,a34769a,a34773a,a34774a,a34777a,a34780a,a34781a,a34782a,a34786a,a34787a,a34790a,a34793a,a34794a,a34795a,a34799a,a34800a,a34803a,a34806a,a34807a,a34808a,a34812a,a34813a,a34816a,a34819a,a34820a,a34821a,a34825a,a34826a,a34829a,a34832a,a34833a,a34834a,a34838a,a34839a,a34842a,a34845a,a34846a,a34847a,a34851a,a34852a,a34855a,a34858a,a34859a,a34860a,a34864a,a34865a,a34868a,a34871a,a34872a,a34873a,a34877a,a34878a,a34881a,a34884a,a34885a,a34886a,a34890a,a34891a,a34894a,a34897a,a34898a,a34899a,a34903a,a34904a,a34907a,a34910a,a34911a,a34912a,a34916a,a34917a,a34920a,a34923a,a34924a,a34925a,a34929a,a34930a,a34933a,a34936a,a34937a,a34938a,a34942a,a34943a,a34946a,a34949a,a34950a,a34951a,a34955a,a34956a,a34959a,a34962a,a34963a,a34964a,a34968a,a34969a,a34972a,a34975a,a34976a,a34977a,a34981a,a34982a,a34985a,a34988a,a34989a,a34990a,a34994a,a34995a,a34998a,a35001a,a35002a,a35003a,a35007a,a35008a,a35011a,a35014a,a35015a,a35016a,a35020a,a35021a,a35024a,a35027a,a35028a,a35029a,a35033a,a35034a,a35037a,a35040a,a35041a,a35042a,a35046a,a35047a,a35050a,a35053a,a35054a,a35055a,a35059a,a35060a,a35063a,a35066a,a35067a,a35068a,a35072a,a35073a,a35076a,a35079a,a35080a,a35081a,a35085a,a35086a,a35089a,a35092a,a35093a,a35094a,a35098a,a35099a,a35102a,a35105a,a35106a,a35107a,a35111a,a35112a,a35115a,a35118a,a35119a,a35120a,a35124a,a35125a,a35128a,a35131a,a35132a,a35133a,a35137a,a35138a,a35141a,a35144a,a35145a,a35146a,a35150a,a35151a,a35154a,a35157a,a35158a,a35159a,a35163a,a35164a,a35167a,a35170a,a35171a,a35172a,a35176a,a35177a,a35180a,a35183a,a35184a,a35185a,a35189a,a35190a,a35193a,a35196a,a35197a,a35198a,a35202a,a35203a,a35206a,a35209a,a35210a,a35211a,a35215a,a35216a,a35219a,a35222a,a35223a,a35224a,a35228a,a35229a,a35232a,a35235a,a35236a,a35237a,a35241a,a35242a,a35245a,a35248a,a35249a,a35250a,a35254a,a35255a,a35258a,a35261a,a35262a,a35263a,a35267a,a35268a,a35271a,a35274a,a35275a,a35276a,a35280a,a35281a,a35284a,a35287a,a35288a,a35289a,a35293a,a35294a,a35297a,a35300a,a35301a,a35302a,a35306a,a35307a,a35310a,a35313a,a35314a,a35315a,a35319a,a35320a,a35323a,a35326a,a35327a,a35328a,a35332a,a35333a,a35336a,a35339a,a35340a,a35341a,a35345a,a35346a,a35349a,a35352a,a35353a,a35354a,a35358a,a35359a,a35362a,a35365a,a35366a,a35367a,a35371a,a35372a,a35375a,a35378a,a35379a,a35380a,a35384a,a35385a,a35388a,a35391a,a35392a,a35393a,a35397a,a35398a,a35401a,a35404a,a35405a,a35406a,a35410a,a35411a,a35414a,a35417a,a35418a,a35419a,a35423a,a35424a,a35427a,a35430a,a35431a,a35432a,a35436a,a35437a,a35440a,a35443a,a35444a,a35445a,a35449a,a35450a,a35453a,a35456a,a35457a,a35458a,a35462a,a35463a,a35466a,a35469a,a35470a,a35471a,a35475a,a35476a,a35479a,a35482a,a35483a,a35484a,a35488a,a35489a,a35492a,a35495a,a35496a,a35497a,a35501a,a35502a,a35505a,a35508a,a35509a,a35510a,a35514a,a35515a,a35518a,a35521a,a35522a,a35523a,a35527a,a35528a,a35531a,a35534a,a35535a,a35536a,a35540a,a35541a,a35544a,a35547a,a35548a,a35549a,a35553a,a35554a,a35557a,a35560a,a35561a,a35562a,a35566a,a35567a,a35570a,a35573a,a35574a,a35575a,a35579a,a35580a,a35583a,a35586a,a35587a,a35588a,a35592a,a35593a,a35596a,a35599a,a35600a,a35601a,a35605a,a35606a,a35609a,a35612a,a35613a,a35614a,a35618a,a35619a,a35622a,a35625a,a35626a,a35627a,a35631a,a35632a,a35635a,a35638a,a35639a,a35640a,a35644a,a35645a,a35648a,a35651a,a35652a,a35653a,a35657a,a35658a,a35661a,a35664a,a35665a,a35666a,a35670a,a35671a,a35674a,a35677a,a35678a,a35679a,a35683a,a35684a,a35687a,a35690a,a35691a,a35692a,a35696a,a35697a,a35700a,a35703a,a35704a,a35705a,a35709a,a35710a,a35713a,a35716a,a35717a,a35718a,a35722a,a35723a,a35726a,a35729a,a35730a,a35731a,a35735a,a35736a,a35739a,a35742a,a35743a,a35744a,a35748a,a35749a,a35752a,a35755a,a35756a,a35757a,a35761a,a35762a,a35765a,a35768a,a35769a,a35770a,a35774a,a35775a,a35778a,a35781a,a35782a,a35783a,a35787a,a35788a,a35791a,a35794a,a35795a,a35796a,a35800a,a35801a,a35804a,a35807a,a35808a,a35809a,a35813a,a35814a,a35817a,a35820a,a35821a,a35822a,a35826a,a35827a,a35830a,a35833a,a35834a,a35835a,a35839a,a35840a,a35843a,a35846a,a35847a,a35848a,a35852a,a35853a,a35856a,a35859a,a35860a,a35861a,a35865a,a35866a,a35869a,a35872a,a35873a,a35874a,a35878a,a35879a,a35882a,a35885a,a35886a,a35887a,a35891a,a35892a,a35895a,a35898a,a35899a,a35900a,a35904a,a35905a,a35908a,a35911a,a35912a,a35913a,a35917a,a35918a,a35921a,a35924a,a35925a,a35926a,a35930a,a35931a,a35934a,a35937a,a35938a,a35939a,a35943a,a35944a,a35947a,a35950a,a35951a,a35952a,a35956a,a35957a,a35960a,a35963a,a35964a,a35965a,a35969a,a35970a,a35973a,a35976a,a35977a,a35978a,a35982a,a35983a,a35986a,a35989a,a35990a,a35991a,a35995a,a35996a,a35999a,a36002a,a36003a,a36004a,a36008a,a36009a,a36012a,a36015a,a36016a,a36017a,a36021a,a36022a,a36025a,a36028a,a36029a,a36030a,a36034a,a36035a,a36038a,a36041a,a36042a,a36043a,a36047a,a36048a,a36051a,a36054a,a36055a,a36056a,a36060a,a36061a,a36064a,a36067a,a36068a,a36069a,a36073a,a36074a,a36077a,a36080a,a36081a,a36082a,a36086a,a36087a,a36090a,a36093a,a36094a,a36095a,a36099a,a36100a,a36103a,a36106a,a36107a,a36108a,a36112a,a36113a,a36116a,a36119a,a36120a,a36121a,a36125a,a36126a,a36129a,a36132a,a36133a,a36134a,a36138a,a36139a,a36142a,a36145a,a36146a,a36147a,a36151a,a36152a,a36155a,a36158a,a36159a,a36160a,a36164a,a36165a,a36168a,a36171a,a36172a,a36173a,a36177a,a36178a,a36181a,a36184a,a36185a,a36186a,a36190a,a36191a,a36194a,a36197a,a36198a,a36199a,a36203a,a36204a,a36207a,a36210a,a36211a,a36212a,a36216a,a36217a,a36220a,a36223a,a36224a,a36225a,a36229a,a36230a,a36233a,a36236a,a36237a,a36238a,a36242a,a36243a,a36246a,a36249a,a36250a,a36251a,a36255a,a36256a,a36259a,a36262a,a36263a,a36264a,a36268a,a36269a,a36272a,a36275a,a36276a,a36277a,a36281a,a36282a,a36285a,a36288a,a36289a,a36290a,a36294a,a36295a,a36298a,a36301a,a36302a,a36303a,a36307a,a36308a,a36311a,a36314a,a36315a,a36316a,a36320a,a36321a,a36324a,a36327a,a36328a,a36329a,a36333a,a36334a,a36337a,a36340a,a36341a,a36342a,a36346a,a36347a,a36350a,a36353a,a36354a,a36355a,a36359a,a36360a,a36363a,a36366a,a36367a,a36368a,a36372a,a36373a,a36376a,a36379a,a36380a,a36381a,a36385a,a36386a,a36389a,a36392a,a36393a,a36394a,a36398a,a36399a,a36402a,a36405a,a36406a,a36407a,a36411a,a36412a,a36415a,a36418a,a36419a,a36420a,a36424a,a36425a,a36428a,a36431a,a36432a,a36433a,a36437a,a36438a,a36441a,a36444a,a36445a,a36446a,a36450a,a36451a,a36454a,a36457a,a36458a,a36459a,a36463a,a36464a,a36467a,a36470a,a36471a,a36472a,a36476a,a36477a,a36480a,a36483a,a36484a,a36485a,a36489a,a36490a,a36493a,a36496a,a36497a,a36498a,a36502a,a36503a,a36506a,a36509a,a36510a,a36511a,a36515a,a36516a,a36519a,a36522a,a36523a,a36524a,a36528a,a36529a,a36532a,a36535a,a36536a,a36537a,a36541a,a36542a,a36545a,a36548a,a36549a,a36550a,a36554a,a36555a,a36558a,a36561a,a36562a,a36563a,a36567a,a36568a,a36571a,a36574a,a36575a,a36576a,a36580a,a36581a,a36584a,a36587a,a36588a,a36589a,a36593a,a36594a,a36597a,a36600a,a36601a,a36602a,a36606a,a36607a,a36610a,a36613a,a36614a,a36615a,a36619a,a36620a,a36623a,a36626a,a36627a,a36628a,a36632a,a36633a,a36636a,a36639a,a36640a,a36641a,a36645a,a36646a,a36649a,a36652a,a36653a,a36654a,a36658a,a36659a,a36662a,a36665a,a36666a,a36667a,a36671a,a36672a,a36675a,a36678a,a36679a,a36680a,a36684a,a36685a,a36688a,a36691a,a36692a,a36693a,a36697a,a36698a,a36701a,a36704a,a36705a,a36706a,a36710a,a36711a,a36714a,a36717a,a36718a,a36719a,a36723a,a36724a,a36727a,a36730a,a36731a,a36732a,a36736a,a36737a,a36740a,a36743a,a36744a,a36745a,a36749a,a36750a,a36753a,a36756a,a36757a,a36758a,a36762a,a36763a,a36766a,a36769a,a36770a,a36771a,a36775a,a36776a,a36779a,a36782a,a36783a,a36784a,a36788a,a36789a,a36792a,a36795a,a36796a,a36797a,a36801a,a36802a,a36805a,a36808a,a36809a,a36810a,a36814a,a36815a,a36818a,a36821a,a36822a,a36823a,a36827a,a36828a,a36831a,a36834a,a36835a,a36836a,a36840a,a36841a,a36844a,a36847a,a36848a,a36849a,a36853a,a36854a,a36857a,a36860a,a36861a,a36862a,a36866a,a36867a,a36870a,a36873a,a36874a,a36875a,a36879a,a36880a,a36883a,a36886a,a36887a,a36888a,a36892a,a36893a,a36896a,a36899a,a36900a,a36901a,a36905a,a36906a,a36909a,a36912a,a36913a,a36914a,a36918a,a36919a,a36922a,a36925a,a36926a,a36927a,a36931a,a36932a,a36935a,a36938a,a36939a,a36940a,a36944a,a36945a,a36948a,a36951a,a36952a,a36953a,a36957a,a36958a,a36961a,a36964a,a36965a,a36966a,a36970a,a36971a,a36974a,a36977a,a36978a,a36979a,a36983a,a36984a,a36987a,a36990a,a36991a,a36992a,a36996a,a36997a,a37000a,a37003a,a37004a,a37005a,a37009a,a37010a,a37013a,a37016a,a37017a,a37018a,a37022a,a37023a,a37026a,a37029a,a37030a,a37031a,a37035a,a37036a,a37039a,a37042a,a37043a,a37044a,a37048a,a37049a,a37052a,a37055a,a37056a,a37057a,a37061a,a37062a,a37065a,a37068a,a37069a,a37070a,a37074a,a37075a,a37078a,a37081a,a37082a,a37083a,a37087a,a37088a,a37091a,a37094a,a37095a,a37096a,a37100a,a37101a,a37104a,a37107a,a37108a,a37109a,a37113a,a37114a,a37117a,a37120a,a37121a,a37122a,a37126a,a37127a,a37130a,a37133a,a37134a,a37135a,a37139a,a37140a,a37143a,a37146a,a37147a,a37148a,a37152a,a37153a,a37156a,a37159a,a37160a,a37161a,a37165a,a37166a,a37169a,a37172a,a37173a,a37174a,a37178a,a37179a,a37182a,a37185a,a37186a,a37187a,a37191a,a37192a,a37195a,a37198a,a37199a,a37200a,a37204a,a37205a,a37208a,a37211a,a37212a,a37213a,a37217a,a37218a,a37221a,a37224a,a37225a,a37226a,a37230a,a37231a,a37234a,a37237a,a37238a,a37239a,a37243a,a37244a,a37247a,a37250a,a37251a,a37252a,a37256a,a37257a,a37260a,a37263a,a37264a,a37265a,a37269a,a37270a,a37273a,a37276a,a37277a,a37278a,a37282a,a37283a,a37286a,a37289a,a37290a,a37291a,a37295a,a37296a,a37299a,a37302a,a37303a,a37304a,a37308a,a37309a,a37312a,a37315a,a37316a,a37317a,a37321a,a37322a,a37325a,a37328a,a37329a,a37330a,a37334a,a37335a,a37338a,a37341a,a37342a,a37343a,a37347a,a37348a,a37351a,a37354a,a37355a,a37356a,a37360a,a37361a,a37364a,a37367a,a37368a,a37369a,a37373a,a37374a,a37377a,a37380a,a37381a,a37382a,a37386a,a37387a,a37390a,a37393a,a37394a,a37395a,a37399a,a37400a,a37403a,a37406a,a37407a,a37408a,a37412a,a37413a,a37416a,a37419a,a37420a,a37421a,a37425a,a37426a,a37429a,a37432a,a37433a,a37434a,a37438a,a37439a,a37442a,a37445a,a37446a,a37447a,a37451a,a37452a,a37455a,a37458a,a37459a,a37460a,a37464a,a37465a,a37468a,a37471a,a37472a,a37473a,a37477a,a37478a,a37481a,a37484a,a37485a,a37486a,a37490a,a37491a,a37494a,a37497a,a37498a,a37499a,a37503a,a37504a,a37507a,a37510a,a37511a,a37512a,a37516a,a37517a,a37520a,a37523a,a37524a,a37525a,a37529a,a37530a,a37533a,a37536a,a37537a,a37538a,a37542a,a37543a,a37546a,a37549a,a37550a,a37551a,a37555a,a37556a,a37559a,a37562a,a37563a,a37564a,a37568a,a37569a,a37572a,a37575a,a37576a,a37577a,a37581a,a37582a,a37585a,a37588a,a37589a,a37590a,a37594a,a37595a,a37598a,a37601a,a37602a,a37603a,a37607a,a37608a,a37611a,a37614a,a37615a,a37616a,a37620a,a37621a,a37624a,a37627a,a37628a,a37629a,a37633a,a37634a,a37637a,a37640a,a37641a,a37642a,a37646a,a37647a,a37650a,a37653a,a37654a,a37655a,a37659a,a37660a,a37663a,a37666a,a37667a,a37668a,a37672a,a37673a,a37676a,a37679a,a37680a,a37681a,a37685a,a37686a,a37689a,a37692a,a37693a,a37694a,a37698a,a37699a,a37702a,a37705a,a37706a,a37707a,a37711a,a37712a,a37715a,a37718a,a37719a,a37720a,a37724a,a37725a,a37728a,a37731a,a37732a,a37733a,a37737a,a37738a,a37741a,a37744a,a37745a,a37746a,a37750a,a37751a,a37754a,a37757a,a37758a,a37759a,a37763a,a37764a,a37767a,a37770a,a37771a,a37772a,a37776a,a37777a,a37780a,a37783a,a37784a,a37785a,a37789a,a37790a,a37793a,a37796a,a37797a,a37798a,a37802a,a37803a,a37806a,a37809a,a37810a,a37811a,a37815a,a37816a,a37819a,a37822a,a37823a,a37824a,a37828a,a37829a,a37832a,a37835a,a37836a,a37837a,a37840a,a37843a,a37844a,a37847a,a37850a,a37851a,a37852a,a37856a,a37857a,a37860a,a37863a,a37864a,a37865a,a37868a,a37871a,a37872a,a37875a,a37878a,a37879a,a37880a,a37884a,a37885a,a37888a,a37891a,a37892a,a37893a,a37896a,a37899a,a37900a,a37903a,a37906a,a37907a,a37908a,a37912a,a37913a,a37916a,a37919a,a37920a,a37921a,a37924a,a37927a,a37928a,a37931a,a37934a,a37935a,a37936a,a37940a,a37941a,a37944a,a37947a,a37948a,a37949a,a37952a,a37955a,a37956a,a37959a,a37962a,a37963a,a37964a,a37968a,a37969a,a37972a,a37975a,a37976a,a37977a,a37980a,a37983a,a37984a,a37987a,a37990a,a37991a,a37992a,a37996a,a37997a,a38000a,a38003a,a38004a,a38005a,a38008a,a38011a,a38012a,a38015a,a38018a,a38019a,a38020a,a38024a,a38025a,a38028a,a38031a,a38032a,a38033a,a38036a,a38039a,a38040a,a38043a,a38046a,a38047a,a38048a,a38052a,a38053a,a38056a,a38059a,a38060a,a38061a,a38064a,a38067a,a38068a,a38071a,a38074a,a38075a,a38076a,a38080a,a38081a,a38084a,a38087a,a38088a,a38089a,a38092a,a38095a,a38096a,a38099a,a38102a,a38103a,a38104a,a38108a,a38109a,a38112a,a38115a,a38116a,a38117a,a38120a,a38123a,a38124a,a38127a,a38130a,a38131a,a38132a,a38136a,a38137a,a38140a,a38143a,a38144a,a38145a,a38148a,a38151a,a38152a,a38155a,a38158a,a38159a,a38160a,a38164a,a38165a,a38168a,a38171a,a38172a,a38173a,a38176a,a38179a,a38180a,a38183a,a38186a,a38187a,a38188a,a38192a,a38193a,a38196a,a38199a,a38200a,a38201a,a38204a,a38207a,a38208a,a38211a,a38214a,a38215a,a38216a,a38220a,a38221a,a38224a,a38227a,a38228a,a38229a,a38232a,a38235a,a38236a,a38239a,a38242a,a38243a,a38244a,a38248a,a38249a,a38252a,a38255a,a38256a,a38257a,a38260a,a38263a,a38264a,a38267a,a38270a,a38271a,a38272a,a38276a,a38277a,a38280a,a38283a,a38284a,a38285a,a38288a,a38291a,a38292a,a38295a,a38298a,a38299a,a38300a,a38304a,a38305a,a38308a,a38311a,a38312a,a38313a,a38316a,a38319a,a38320a,a38323a,a38326a,a38327a,a38328a,a38332a,a38333a,a38336a,a38339a,a38340a,a38341a,a38344a,a38347a,a38348a,a38351a,a38354a,a38355a,a38356a,a38360a,a38361a,a38364a,a38367a,a38368a,a38369a,a38372a,a38375a,a38376a,a38379a,a38382a,a38383a,a38384a,a38388a,a38389a,a38392a,a38395a,a38396a,a38397a,a38400a,a38403a,a38404a,a38407a,a38410a,a38411a,a38412a,a38416a,a38417a,a38420a,a38423a,a38424a,a38425a,a38428a,a38431a,a38432a,a38435a,a38438a,a38439a,a38440a,a38444a,a38445a,a38448a,a38451a,a38452a,a38453a,a38456a,a38459a,a38460a,a38463a,a38466a,a38467a,a38468a,a38472a,a38473a,a38476a,a38479a,a38480a,a38481a,a38484a,a38487a,a38488a,a38491a,a38494a,a38495a,a38496a,a38500a,a38501a,a38504a,a38507a,a38508a,a38509a,a38512a,a38515a,a38516a,a38519a,a38522a,a38523a,a38524a,a38528a,a38529a,a38532a,a38535a,a38536a,a38537a,a38540a,a38543a,a38544a,a38547a,a38550a,a38551a,a38552a,a38556a,a38557a,a38560a,a38563a,a38564a,a38565a,a38568a,a38571a,a38572a,a38575a,a38578a,a38579a,a38580a,a38584a,a38585a,a38588a,a38591a,a38592a,a38593a,a38596a,a38599a,a38600a,a38603a,a38606a,a38607a,a38608a,a38612a,a38613a,a38616a,a38619a,a38620a,a38621a,a38624a,a38627a,a38628a,a38631a,a38634a,a38635a,a38636a,a38640a,a38641a,a38644a,a38647a,a38648a,a38649a,a38652a,a38655a,a38656a,a38659a,a38662a,a38663a,a38664a,a38668a,a38669a,a38672a,a38675a,a38676a,a38677a,a38680a,a38683a,a38684a,a38687a,a38690a,a38691a,a38692a,a38696a,a38697a,a38700a,a38703a,a38704a,a38705a,a38708a,a38711a,a38712a,a38715a,a38718a,a38719a,a38720a,a38724a,a38725a,a38728a,a38731a,a38732a,a38733a,a38736a,a38739a,a38740a,a38743a,a38746a,a38747a,a38748a,a38752a,a38753a,a38756a,a38759a,a38760a,a38761a,a38764a,a38767a,a38768a,a38771a,a38774a,a38775a,a38776a,a38780a,a38781a,a38784a,a38787a,a38788a,a38789a,a38792a,a38795a,a38796a,a38799a,a38802a,a38803a,a38804a,a38808a,a38809a,a38812a,a38815a,a38816a,a38817a,a38820a,a38823a,a38824a,a38827a,a38830a,a38831a,a38832a,a38836a,a38837a,a38840a,a38843a,a38844a,a38845a,a38848a,a38851a,a38852a,a38855a,a38858a,a38859a,a38860a,a38864a,a38865a,a38868a,a38871a,a38872a,a38873a,a38876a,a38879a,a38880a,a38883a,a38886a,a38887a,a38888a,a38892a,a38893a,a38896a,a38899a,a38900a,a38901a,a38904a,a38907a,a38908a,a38911a,a38914a,a38915a,a38916a,a38920a,a38921a,a38924a,a38927a,a38928a,a38929a,a38932a,a38935a,a38936a,a38939a,a38942a,a38943a,a38944a,a38948a,a38949a,a38952a,a38955a,a38956a,a38957a,a38960a,a38963a,a38964a,a38967a,a38970a,a38971a,a38972a,a38976a,a38977a,a38980a,a38983a,a38984a,a38985a,a38988a,a38991a,a38992a,a38995a,a38998a,a38999a,a39000a,a39004a,a39005a,a39008a,a39011a,a39012a,a39013a,a39016a,a39019a,a39020a,a39023a,a39026a,a39027a,a39028a,a39032a,a39033a,a39036a,a39039a,a39040a,a39041a,a39044a,a39047a,a39048a,a39051a,a39054a,a39055a,a39056a,a39060a,a39061a,a39064a,a39067a,a39068a,a39069a,a39072a,a39075a,a39076a,a39079a,a39082a,a39083a,a39084a,a39088a,a39089a,a39092a,a39095a,a39096a,a39097a,a39100a,a39103a,a39104a,a39107a,a39110a,a39111a,a39112a,a39116a,a39117a,a39120a,a39123a,a39124a,a39125a,a39128a,a39131a,a39132a,a39135a,a39138a,a39139a,a39140a,a39144a,a39145a,a39148a,a39151a,a39152a,a39153a,a39156a,a39159a,a39160a,a39163a,a39166a,a39167a,a39168a,a39172a,a39173a,a39176a,a39179a,a39180a,a39181a,a39184a,a39187a,a39188a,a39191a,a39194a,a39195a,a39196a,a39200a,a39201a,a39204a,a39207a,a39208a,a39209a,a39212a,a39215a,a39216a,a39219a,a39222a,a39223a,a39224a,a39228a,a39229a,a39232a,a39235a,a39236a,a39237a,a39240a,a39243a,a39244a,a39247a,a39250a,a39251a,a39252a,a39256a,a39257a,a39260a,a39263a,a39264a,a39265a,a39268a,a39271a,a39272a,a39275a,a39278a,a39279a,a39280a,a39284a,a39285a,a39288a,a39291a,a39292a,a39293a,a39296a,a39299a,a39300a,a39303a,a39306a,a39307a,a39308a,a39312a,a39313a,a39316a,a39319a,a39320a,a39321a,a39324a,a39327a,a39328a,a39331a,a39334a,a39335a,a39336a,a39340a,a39341a,a39344a,a39347a,a39348a,a39349a,a39352a,a39355a,a39356a,a39359a,a39362a,a39363a,a39364a,a39368a,a39369a,a39372a,a39375a,a39376a,a39377a,a39380a,a39383a,a39384a,a39387a,a39390a,a39391a,a39392a,a39396a,a39397a,a39400a,a39403a,a39404a,a39405a,a39408a,a39411a,a39412a,a39415a,a39418a,a39419a,a39420a,a39424a,a39425a,a39428a,a39431a,a39432a,a39433a,a39436a,a39439a,a39440a,a39443a,a39446a,a39447a,a39448a,a39452a,a39453a,a39456a,a39459a,a39460a,a39461a,a39464a,a39467a,a39468a,a39471a,a39474a,a39475a,a39476a,a39480a,a39481a,a39484a,a39487a,a39488a,a39489a,a39492a,a39495a,a39496a,a39499a,a39502a,a39503a,a39504a,a39508a,a39509a,a39512a,a39515a,a39516a,a39517a,a39520a,a39523a,a39524a,a39527a,a39530a,a39531a,a39532a,a39536a,a39537a,a39540a,a39543a,a39544a,a39545a,a39548a,a39551a,a39552a,a39555a,a39558a,a39559a,a39560a,a39564a,a39565a,a39568a,a39571a,a39572a,a39573a,a39576a,a39579a,a39580a,a39583a,a39586a,a39587a,a39588a,a39592a,a39593a,a39596a,a39599a,a39600a,a39601a,a39604a,a39607a,a39608a,a39611a,a39614a,a39615a,a39616a,a39620a,a39621a,a39624a,a39627a,a39628a,a39629a,a39632a,a39635a,a39636a,a39639a,a39642a,a39643a,a39644a,a39648a,a39649a,a39652a,a39655a,a39656a,a39657a,a39660a,a39663a,a39664a,a39667a,a39670a,a39671a,a39672a,a39676a,a39677a,a39680a,a39683a,a39684a,a39685a,a39688a,a39691a,a39692a,a39695a,a39698a,a39699a,a39700a,a39704a,a39705a,a39708a,a39711a,a39712a,a39713a,a39716a,a39719a,a39720a,a39723a,a39726a,a39727a,a39728a,a39732a,a39733a,a39736a,a39739a,a39740a,a39741a,a39744a,a39747a,a39748a,a39751a,a39754a,a39755a,a39756a,a39760a,a39761a,a39764a,a39767a,a39768a,a39769a,a39772a,a39775a,a39776a,a39779a,a39782a,a39783a,a39784a,a39788a,a39789a,a39792a,a39795a,a39796a,a39797a,a39800a,a39803a,a39804a,a39807a,a39810a,a39811a,a39812a,a39816a,a39817a,a39820a,a39823a,a39824a,a39825a,a39828a,a39831a,a39832a,a39835a,a39838a,a39839a,a39840a,a39844a,a39845a,a39848a,a39851a,a39852a,a39853a,a39856a,a39859a,a39860a,a39863a,a39866a,a39867a,a39868a,a39872a,a39873a,a39876a,a39879a,a39880a,a39881a,a39884a,a39887a,a39888a,a39891a,a39894a,a39895a,a39896a,a39900a,a39901a,a39904a,a39907a,a39908a,a39909a,a39912a,a39915a,a39916a,a39919a,a39922a,a39923a,a39924a,a39928a,a39929a,a39932a,a39935a,a39936a,a39937a,a39940a,a39943a,a39944a,a39947a,a39950a,a39951a,a39952a,a39956a,a39957a,a39960a,a39963a,a39964a,a39965a,a39968a,a39971a,a39972a,a39975a,a39978a,a39979a,a39980a,a39984a,a39985a,a39988a,a39991a,a39992a,a39993a,a39996a,a39999a,a40000a,a40003a,a40006a,a40007a,a40008a,a40012a,a40013a,a40016a,a40019a,a40020a,a40021a,a40024a,a40027a,a40028a,a40031a,a40034a,a40035a,a40036a,a40040a,a40041a,a40044a,a40047a,a40048a,a40049a,a40052a,a40055a,a40056a,a40059a,a40062a,a40063a,a40064a,a40068a,a40069a,a40072a,a40075a,a40076a,a40077a,a40080a,a40083a,a40084a,a40087a,a40090a,a40091a,a40092a,a40096a,a40097a,a40100a,a40103a,a40104a,a40105a,a40108a,a40111a,a40112a,a40115a,a40118a,a40119a,a40120a,a40124a,a40125a,a40128a,a40131a,a40132a,a40133a,a40136a,a40139a,a40140a,a40143a,a40146a,a40147a,a40148a,a40152a,a40153a,a40156a,a40159a,a40160a,a40161a,a40164a,a40167a,a40168a,a40171a,a40174a,a40175a,a40176a,a40180a,a40181a,a40184a,a40187a,a40188a,a40189a,a40192a,a40195a,a40196a,a40199a,a40202a,a40203a,a40204a,a40208a,a40209a,a40212a,a40215a,a40216a,a40217a,a40220a,a40223a,a40224a,a40227a,a40230a,a40231a,a40232a,a40236a,a40237a,a40240a,a40243a,a40244a,a40245a,a40248a,a40251a,a40252a,a40255a,a40258a,a40259a,a40260a,a40264a,a40265a,a40268a,a40271a,a40272a,a40273a,a40276a,a40279a,a40280a,a40283a,a40286a,a40287a,a40288a,a40292a,a40293a,a40296a,a40299a,a40300a,a40301a,a40304a,a40307a,a40308a,a40311a,a40314a,a40315a,a40316a,a40320a,a40321a,a40324a,a40327a,a40328a,a40329a,a40332a,a40335a,a40336a,a40339a,a40342a,a40343a,a40344a,a40348a,a40349a,a40352a,a40355a,a40356a,a40357a,a40360a,a40363a,a40364a,a40367a,a40370a,a40371a,a40372a,a40376a,a40377a,a40380a,a40383a,a40384a,a40385a,a40388a,a40391a,a40392a,a40395a,a40398a,a40399a,a40400a,a40404a,a40405a,a40408a,a40411a,a40412a,a40413a,a40416a,a40419a,a40420a,a40423a,a40426a,a40427a,a40428a,a40432a,a40433a,a40436a,a40439a,a40440a,a40441a,a40444a,a40447a,a40448a,a40451a,a40454a,a40455a,a40456a,a40460a,a40461a,a40464a,a40467a,a40468a,a40469a,a40472a,a40475a,a40476a,a40479a,a40482a,a40483a,a40484a,a40488a,a40489a,a40492a,a40495a,a40496a,a40497a,a40500a,a40503a,a40504a,a40507a,a40510a,a40511a,a40512a,a40516a,a40517a,a40520a,a40523a,a40524a,a40525a,a40528a,a40531a,a40532a,a40535a,a40538a,a40539a,a40540a,a40544a,a40545a,a40548a,a40551a,a40552a,a40553a,a40556a,a40559a,a40560a,a40563a,a40566a,a40567a,a40568a,a40572a,a40573a,a40576a,a40579a,a40580a,a40581a,a40584a,a40587a,a40588a,a40591a,a40594a,a40595a,a40596a,a40600a,a40601a,a40604a,a40607a,a40608a,a40609a,a40612a,a40615a,a40616a,a40619a,a40622a,a40623a,a40624a,a40628a,a40629a,a40632a,a40635a,a40636a,a40637a,a40640a,a40643a,a40644a,a40647a,a40650a,a40651a,a40652a,a40656a,a40657a,a40660a,a40663a,a40664a,a40665a,a40668a,a40671a,a40672a,a40675a,a40678a,a40679a,a40680a,a40684a,a40685a,a40688a,a40691a,a40692a,a40693a,a40696a,a40699a,a40700a,a40703a,a40706a,a40707a,a40708a,a40712a,a40713a,a40716a,a40719a,a40720a,a40721a,a40724a,a40727a,a40728a,a40731a,a40734a,a40735a,a40736a,a40740a,a40741a,a40744a,a40747a,a40748a,a40749a,a40752a,a40755a,a40756a,a40759a,a40762a,a40763a,a40764a,a40768a,a40769a,a40772a,a40775a,a40776a,a40777a,a40780a,a40783a,a40784a,a40787a,a40790a,a40791a,a40792a,a40796a,a40797a,a40800a,a40803a,a40804a,a40805a,a40808a,a40811a,a40812a,a40815a,a40818a,a40819a,a40820a,a40824a,a40825a,a40828a,a40831a,a40832a,a40833a,a40836a,a40839a,a40840a,a40843a,a40846a,a40847a,a40848a,a40852a,a40853a,a40856a,a40859a,a40860a,a40861a,a40864a,a40867a,a40868a,a40871a,a40874a,a40875a,a40876a,a40880a,a40881a,a40884a,a40887a,a40888a,a40889a,a40892a,a40895a,a40896a,a40899a,a40902a,a40903a,a40904a,a40908a,a40909a,a40912a,a40915a,a40916a,a40917a,a40920a,a40923a,a40924a,a40927a,a40930a,a40931a,a40932a,a40936a,a40937a,a40940a,a40943a,a40944a,a40945a,a40948a,a40951a,a40952a,a40955a,a40958a,a40959a,a40960a,a40964a,a40965a,a40968a,a40971a,a40972a,a40973a,a40976a,a40979a,a40980a,a40983a,a40986a,a40987a,a40988a,a40992a,a40993a,a40996a,a40999a,a41000a,a41001a,a41004a,a41007a,a41008a,a41011a,a41014a,a41015a,a41016a,a41020a,a41021a,a41024a,a41027a,a41028a,a41029a,a41032a,a41035a,a41036a,a41039a,a41042a,a41043a,a41044a,a41048a,a41049a,a41052a,a41055a,a41056a,a41057a,a41060a,a41063a,a41064a,a41067a,a41070a,a41071a,a41072a,a41076a,a41077a,a41080a,a41083a,a41084a,a41085a,a41088a,a41091a,a41092a,a41095a,a41098a,a41099a,a41100a,a41104a,a41105a,a41108a,a41111a,a41112a,a41113a,a41116a,a41119a,a41120a,a41123a,a41126a,a41127a,a41128a,a41132a,a41133a,a41136a,a41139a,a41140a,a41141a,a41144a,a41147a,a41148a,a41151a,a41154a,a41155a,a41156a,a41160a,a41161a,a41164a,a41167a,a41168a,a41169a,a41172a,a41175a,a41176a,a41179a,a41182a,a41183a,a41184a,a41188a,a41189a,a41192a,a41195a,a41196a,a41197a,a41200a,a41203a,a41204a,a41207a,a41210a,a41211a,a41212a,a41216a,a41217a,a41220a,a41223a,a41224a,a41225a,a41228a,a41231a,a41232a,a41235a,a41238a,a41239a,a41240a,a41244a,a41245a,a41248a,a41251a,a41252a,a41253a,a41256a,a41259a,a41260a,a41263a,a41266a,a41267a,a41268a,a41272a,a41273a,a41276a,a41279a,a41280a,a41281a,a41284a,a41287a,a41288a,a41291a,a41294a,a41295a,a41296a,a41300a,a41301a,a41304a,a41307a,a41308a,a41309a,a41312a,a41315a,a41316a,a41319a,a41322a,a41323a,a41324a,a41328a,a41329a,a41332a,a41335a,a41336a,a41337a,a41340a,a41343a,a41344a,a41347a,a41350a,a41351a,a41352a,a41356a,a41357a,a41360a,a41363a,a41364a,a41365a,a41368a,a41371a,a41372a,a41375a,a41378a,a41379a,a41380a,a41384a,a41385a,a41388a,a41391a,a41392a,a41393a,a41396a,a41399a,a41400a,a41403a,a41406a,a41407a,a41408a,a41412a,a41413a,a41416a,a41419a,a41420a,a41421a,a41424a,a41427a,a41428a,a41431a,a41434a,a41435a,a41436a,a41440a,a41441a,a41444a,a41447a,a41448a,a41449a,a41452a,a41455a,a41456a,a41459a,a41462a,a41463a,a41464a,a41468a,a41469a,a41472a,a41475a,a41476a,a41477a,a41480a,a41483a,a41484a,a41487a,a41490a,a41491a,a41492a,a41496a,a41497a,a41500a,a41503a,a41504a,a41505a,a41508a,a41511a,a41512a,a41515a,a41518a,a41519a,a41520a,a41524a,a41525a,a41528a,a41531a,a41532a,a41533a,a41536a,a41539a,a41540a,a41543a,a41546a,a41547a,a41548a,a41552a,a41553a,a41556a,a41559a,a41560a,a41561a,a41564a,a41567a,a41568a,a41571a,a41574a,a41575a,a41576a,a41580a,a41581a,a41584a,a41587a,a41588a,a41589a,a41592a,a41595a,a41596a,a41599a,a41602a,a41603a,a41604a,a41608a,a41609a,a41612a,a41615a,a41616a,a41617a,a41620a,a41623a,a41624a,a41627a,a41630a,a41631a,a41632a,a41636a,a41637a,a41640a,a41643a,a41644a,a41645a,a41648a,a41651a,a41652a,a41655a,a41658a,a41659a,a41660a,a41664a,a41665a,a41668a,a41671a,a41672a,a41673a,a41676a,a41679a,a41680a,a41683a,a41686a,a41687a,a41688a,a41692a,a41693a,a41696a,a41699a,a41700a,a41701a,a41704a,a41707a,a41708a,a41711a,a41714a,a41715a,a41716a,a41720a,a41721a,a41724a,a41727a,a41728a,a41729a,a41732a,a41735a,a41736a,a41739a,a41742a,a41743a,a41744a,a41748a,a41749a,a41752a,a41755a,a41756a,a41757a,a41760a,a41763a,a41764a,a41767a,a41770a,a41771a,a41772a,a41776a,a41777a,a41780a,a41783a,a41784a,a41785a,a41788a,a41791a,a41792a,a41795a,a41798a,a41799a,a41800a,a41804a,a41805a,a41808a,a41811a,a41812a,a41813a,a41816a,a41819a,a41820a,a41823a,a41826a,a41827a,a41828a,a41832a,a41833a,a41836a,a41839a,a41840a,a41841a,a41844a,a41847a,a41848a,a41851a,a41854a,a41855a,a41856a,a41860a,a41861a,a41864a,a41867a,a41868a,a41869a,a41872a,a41875a,a41876a,a41879a,a41882a,a41883a,a41884a,a41888a,a41889a,a41892a,a41895a,a41896a,a41897a,a41900a,a41903a,a41904a,a41907a,a41910a,a41911a,a41912a,a41916a,a41917a,a41920a,a41923a,a41924a,a41925a,a41928a,a41931a,a41932a,a41935a,a41938a,a41939a,a41940a,a41944a,a41945a,a41948a,a41951a,a41952a,a41953a,a41956a,a41959a,a41960a,a41963a,a41966a,a41967a,a41968a,a41972a,a41973a,a41976a,a41979a,a41980a,a41981a,a41984a,a41987a,a41988a,a41991a,a41994a,a41995a,a41996a,a42000a,a42001a,a42004a,a42007a,a42008a,a42009a,a42012a,a42015a,a42016a,a42019a,a42022a,a42023a,a42024a,a42028a,a42029a,a42032a,a42035a,a42036a,a42037a,a42040a,a42043a,a42044a,a42047a,a42050a,a42051a,a42052a,a42056a,a42057a,a42060a,a42063a,a42064a,a42065a,a42068a,a42071a,a42072a,a42075a,a42078a,a42079a,a42080a,a42084a,a42085a,a42088a,a42091a,a42092a,a42093a,a42096a,a42099a,a42100a,a42103a,a42106a,a42107a,a42108a,a42112a,a42113a,a42116a,a42119a,a42120a,a42121a,a42124a,a42127a,a42128a,a42131a,a42134a,a42135a,a42136a,a42140a,a42141a,a42144a,a42147a,a42148a,a42149a,a42152a,a42155a,a42156a,a42159a,a42162a,a42163a,a42164a,a42168a,a42169a,a42172a,a42175a,a42176a,a42177a,a42180a,a42183a,a42184a,a42187a,a42190a,a42191a,a42192a,a42196a,a42197a,a42200a,a42203a,a42204a,a42205a,a42208a,a42211a,a42212a,a42215a,a42218a,a42219a,a42220a,a42224a,a42225a,a42228a,a42231a,a42232a,a42233a,a42236a,a42239a,a42240a,a42243a,a42246a,a42247a,a42248a,a42252a,a42253a,a42256a,a42259a,a42260a,a42261a,a42264a,a42267a,a42268a,a42271a,a42274a,a42275a,a42276a,a42280a,a42281a,a42284a,a42287a,a42288a,a42289a,a42292a,a42295a,a42296a,a42299a,a42302a,a42303a,a42304a,a42308a,a42309a,a42312a,a42315a,a42316a,a42317a,a42320a,a42323a,a42324a,a42327a,a42330a,a42331a,a42332a,a42336a,a42337a,a42340a,a42343a,a42344a,a42345a,a42348a,a42351a,a42352a,a42355a,a42358a,a42359a,a42360a,a42364a,a42365a,a42368a,a42371a,a42372a,a42373a,a42376a,a42379a,a42380a,a42383a,a42386a,a42387a,a42388a,a42392a,a42393a,a42396a,a42399a,a42400a,a42401a,a42404a,a42407a,a42408a,a42411a,a42414a,a42415a,a42416a,a42420a,a42421a,a42424a,a42427a,a42428a,a42429a,a42432a,a42435a,a42436a,a42439a,a42442a,a42443a,a42444a,a42448a,a42449a,a42452a,a42455a,a42456a,a42457a,a42460a,a42463a,a42464a,a42467a,a42470a,a42471a,a42472a,a42476a,a42477a,a42480a,a42483a,a42484a,a42485a,a42488a,a42491a,a42492a,a42495a,a42498a,a42499a,a42500a,a42504a,a42505a,a42508a,a42511a,a42512a,a42513a,a42516a,a42519a,a42520a,a42523a,a42526a,a42527a,a42528a,a42532a,a42533a,a42536a,a42539a,a42540a,a42541a,a42544a,a42547a,a42548a,a42551a,a42554a,a42555a,a42556a,a42560a,a42561a,a42564a,a42567a,a42568a,a42569a,a42572a,a42575a,a42576a,a42579a,a42582a,a42583a,a42584a,a42588a,a42589a,a42592a,a42595a,a42596a,a42597a,a42600a,a42603a,a42604a,a42607a,a42610a,a42611a,a42612a,a42616a,a42617a,a42620a,a42623a,a42624a,a42625a,a42628a,a42631a,a42632a,a42635a,a42638a,a42639a,a42640a,a42644a,a42645a,a42648a,a42651a,a42652a,a42653a,a42656a,a42659a,a42660a,a42663a,a42666a,a42667a,a42668a,a42672a,a42673a,a42676a,a42679a,a42680a,a42681a,a42684a,a42687a,a42688a,a42691a,a42694a,a42695a,a42696a,a42700a,a42701a,a42704a,a42707a,a42708a,a42709a,a42712a,a42715a,a42716a,a42719a,a42722a,a42723a,a42724a,a42728a,a42729a,a42732a,a42735a,a42736a,a42737a,a42740a,a42743a,a42744a,a42747a,a42750a,a42751a,a42752a,a42756a,a42757a,a42760a,a42763a,a42764a,a42765a,a42768a,a42771a,a42772a,a42775a,a42778a,a42779a,a42780a,a42784a,a42785a,a42788a,a42791a,a42792a,a42793a,a42796a,a42799a,a42800a,a42803a,a42806a,a42807a,a42808a,a42812a,a42813a,a42816a,a42819a,a42820a,a42821a,a42824a,a42827a,a42828a,a42831a,a42834a,a42835a,a42836a,a42840a,a42841a,a42844a,a42847a,a42848a,a42849a,a42852a,a42855a,a42856a,a42859a,a42862a,a42863a,a42864a,a42868a,a42869a,a42872a,a42875a,a42876a,a42877a,a42880a,a42883a,a42884a,a42887a,a42890a,a42891a,a42892a,a42896a,a42897a,a42900a,a42903a,a42904a,a42905a,a42908a,a42911a,a42912a,a42915a,a42918a,a42919a,a42920a,a42924a,a42925a,a42928a,a42931a,a42932a,a42933a,a42936a,a42939a,a42940a,a42943a,a42946a,a42947a,a42948a,a42952a,a42953a,a42956a,a42959a,a42960a,a42961a,a42964a,a42967a,a42968a,a42971a,a42974a,a42975a,a42976a,a42980a,a42981a,a42984a,a42987a,a42988a,a42989a,a42992a,a42995a,a42996a,a42999a,a43002a,a43003a,a43004a,a43008a,a43009a,a43012a,a43015a,a43016a,a43017a,a43020a,a43023a,a43024a,a43027a,a43030a,a43031a,a43032a,a43036a,a43037a,a43040a,a43043a,a43044a,a43045a,a43048a,a43051a,a43052a,a43055a,a43058a,a43059a,a43060a,a43064a,a43065a,a43068a,a43071a,a43072a,a43073a,a43076a,a43079a,a43080a,a43083a,a43086a,a43087a,a43088a,a43092a,a43093a,a43096a,a43099a,a43100a,a43101a,a43104a,a43107a,a43108a,a43111a,a43114a,a43115a,a43116a,a43120a,a43121a,a43124a,a43127a,a43128a,a43129a,a43132a,a43135a,a43136a,a43139a,a43142a,a43143a,a43144a,a43148a,a43149a,a43152a,a43155a,a43156a,a43157a,a43160a,a43163a,a43164a,a43167a,a43170a,a43171a,a43172a,a43176a,a43177a,a43180a,a43183a,a43184a,a43185a,a43188a,a43191a,a43192a,a43195a,a43198a,a43199a,a43200a,a43204a,a43205a,a43208a,a43211a,a43212a,a43213a,a43216a,a43219a,a43220a,a43223a,a43226a,a43227a,a43228a,a43232a,a43233a,a43236a,a43239a,a43240a,a43241a,a43244a,a43247a,a43248a,a43251a,a43254a,a43255a,a43256a,a43260a,a43261a,a43264a,a43267a,a43268a,a43269a,a43272a,a43275a,a43276a,a43279a,a43282a,a43283a,a43284a,a43288a,a43289a,a43292a,a43295a,a43296a,a43297a,a43300a,a43303a,a43304a,a43307a,a43310a,a43311a,a43312a,a43316a,a43317a,a43320a,a43323a,a43324a,a43325a,a43328a,a43331a,a43332a,a43335a,a43338a,a43339a,a43340a,a43344a,a43345a,a43348a,a43351a,a43352a,a43353a,a43356a,a43359a,a43360a,a43363a,a43366a,a43367a,a43368a,a43372a,a43373a,a43376a,a43379a,a43380a,a43381a,a43384a,a43387a,a43388a,a43391a,a43394a,a43395a,a43396a,a43400a,a43401a,a43404a,a43407a,a43408a,a43409a,a43412a,a43415a,a43416a,a43419a,a43422a,a43423a,a43424a,a43428a,a43429a,a43432a,a43435a,a43436a,a43437a,a43440a,a43443a,a43444a,a43447a,a43450a,a43451a,a43452a,a43456a,a43457a,a43460a,a43463a,a43464a,a43465a,a43468a,a43471a,a43472a,a43475a,a43478a,a43479a,a43480a,a43484a,a43485a,a43488a,a43491a,a43492a,a43493a,a43496a,a43499a,a43500a,a43503a,a43506a,a43507a,a43508a,a43512a,a43513a,a43516a,a43519a,a43520a,a43521a,a43524a,a43527a,a43528a,a43531a,a43534a,a43535a,a43536a,a43540a,a43541a,a43544a,a43547a,a43548a,a43549a,a43552a,a43555a,a43556a,a43559a,a43562a,a43563a,a43564a,a43568a,a43569a,a43572a,a43575a,a43576a,a43577a,a43580a,a43583a,a43584a,a43587a,a43590a,a43591a,a43592a,a43596a,a43597a,a43600a,a43603a,a43604a,a43605a,a43608a,a43611a,a43612a,a43615a,a43618a,a43619a,a43620a,a43624a,a43625a,a43628a,a43631a,a43632a,a43633a,a43636a,a43639a,a43640a,a43643a,a43646a,a43647a,a43648a,a43652a,a43653a,a43656a,a43659a,a43660a,a43661a,a43664a,a43667a,a43668a,a43671a,a43674a,a43675a,a43676a,a43680a,a43681a,a43684a,a43687a,a43688a,a43689a,a43692a,a43695a,a43696a,a43699a,a43702a,a43703a,a43704a,a43708a,a43709a,a43712a,a43715a,a43716a,a43717a,a43720a,a43723a,a43724a,a43727a,a43730a,a43731a,a43732a,a43736a,a43737a,a43740a,a43743a,a43744a,a43745a,a43748a,a43751a,a43752a,a43755a,a43758a,a43759a,a43760a,a43764a,a43765a,a43768a,a43771a,a43772a,a43773a,a43776a,a43779a,a43780a,a43783a,a43786a,a43787a,a43788a,a43792a,a43793a,a43796a,a43799a,a43800a,a43801a,a43804a,a43807a,a43808a,a43811a,a43814a,a43815a,a43816a,a43820a,a43821a,a43824a,a43827a,a43828a,a43829a,a43832a,a43835a,a43836a,a43839a,a43842a,a43843a,a43844a,a43848a,a43849a,a43852a,a43855a,a43856a,a43857a,a43860a,a43863a,a43864a,a43867a,a43870a,a43871a,a43872a,a43876a,a43877a,a43880a,a43883a,a43884a,a43885a,a43888a,a43891a,a43892a,a43895a,a43898a,a43899a,a43900a,a43904a,a43905a,a43908a,a43911a,a43912a,a43913a,a43916a,a43919a,a43920a,a43923a,a43926a,a43927a,a43928a,a43932a,a43933a,a43936a,a43939a,a43940a,a43941a,a43944a,a43947a,a43948a,a43951a,a43954a,a43955a,a43956a,a43960a,a43961a,a43964a,a43967a,a43968a,a43969a,a43972a,a43975a,a43976a,a43979a,a43982a,a43983a,a43984a,a43988a,a43989a,a43992a,a43995a,a43996a,a43997a,a44000a,a44003a,a44004a,a44007a,a44010a,a44011a,a44012a,a44016a,a44017a,a44020a,a44023a,a44024a,a44025a,a44028a,a44031a,a44032a,a44035a,a44038a,a44039a,a44040a,a44044a,a44045a,a44048a,a44051a,a44052a,a44053a,a44056a,a44059a,a44060a,a44063a,a44066a,a44067a,a44068a,a44072a,a44073a,a44076a,a44079a,a44080a,a44081a,a44084a,a44087a,a44088a,a44091a,a44094a,a44095a,a44096a,a44100a,a44101a,a44104a,a44107a,a44108a,a44109a,a44112a,a44115a,a44116a,a44119a,a44122a,a44123a,a44124a,a44128a,a44129a,a44132a,a44135a,a44136a,a44137a,a44140a,a44143a,a44144a,a44147a,a44150a,a44151a,a44152a,a44156a,a44157a,a44160a,a44163a,a44164a,a44165a,a44168a,a44171a,a44172a,a44175a,a44178a,a44179a,a44180a,a44184a,a44185a,a44188a,a44191a,a44192a,a44193a,a44196a,a44199a,a44200a,a44203a,a44206a,a44207a,a44208a,a44212a,a44213a,a44216a,a44219a,a44220a,a44221a,a44224a,a44227a,a44228a,a44231a,a44234a,a44235a,a44236a,a44240a,a44241a,a44244a,a44247a,a44248a,a44249a,a44252a,a44255a,a44256a,a44259a,a44262a,a44263a,a44264a,a44268a,a44269a,a44272a,a44275a,a44276a,a44277a,a44280a,a44283a,a44284a,a44287a,a44290a,a44291a,a44292a,a44296a,a44297a,a44300a,a44303a,a44304a,a44305a,a44308a,a44311a,a44312a,a44315a,a44318a,a44319a,a44320a,a44324a,a44325a,a44328a,a44331a,a44332a,a44333a,a44336a,a44339a,a44340a,a44343a,a44346a,a44347a,a44348a,a44352a,a44353a,a44356a,a44359a,a44360a,a44361a,a44364a,a44367a,a44368a,a44371a,a44374a,a44375a,a44376a,a44380a,a44381a,a44384a,a44387a,a44388a,a44389a,a44392a,a44395a,a44396a,a44399a,a44402a,a44403a,a44404a,a44408a,a44409a,a44412a,a44415a,a44416a,a44417a,a44420a,a44423a,a44424a,a44427a,a44430a,a44431a,a44432a,a44436a,a44437a,a44440a,a44443a,a44444a,a44445a,a44448a,a44451a,a44452a,a44455a,a44458a,a44459a,a44460a,a44464a,a44465a,a44468a,a44471a,a44472a,a44473a,a44476a,a44479a,a44480a,a44483a,a44486a,a44487a,a44488a,a44492a,a44493a,a44496a,a44499a,a44500a,a44501a,a44504a,a44507a,a44508a,a44511a,a44514a,a44515a,a44516a,a44520a,a44521a,a44524a,a44527a,a44528a,a44529a,a44532a,a44535a,a44536a,a44539a,a44542a,a44543a,a44544a,a44547a,a44550a,a44551a,a44554a,a44557a,a44558a,a44559a,a44562a,a44565a,a44566a,a44569a,a44572a,a44573a,a44574a,a44577a,a44580a,a44581a,a44584a,a44587a,a44588a,a44589a,a44592a,a44595a,a44596a,a44599a,a44602a,a44603a,a44604a,a44607a,a44610a,a44611a,a44614a,a44617a,a44618a,a44619a,a44622a,a44625a,a44626a,a44629a,a44632a,a44633a,a44634a,a44637a,a44640a,a44641a,a44644a,a44647a,a44648a,a44649a,a44652a,a44655a,a44656a,a44659a,a44662a,a44663a,a44664a,a44667a,a44670a,a44671a,a44674a,a44677a,a44678a,a44679a,a44682a,a44685a,a44686a,a44689a,a44692a,a44693a,a44694a,a44697a,a44700a,a44701a,a44704a,a44707a,a44708a,a44709a,a44712a,a44715a,a44716a,a44719a,a44722a,a44723a,a44724a,a44727a,a44730a,a44731a,a44734a,a44737a,a44738a,a44739a,a44742a,a44745a,a44746a,a44749a,a44752a,a44753a,a44754a,a44757a,a44760a,a44761a,a44764a,a44767a,a44768a,a44769a,a44772a,a44775a,a44776a,a44779a,a44782a,a44783a,a44784a,a44787a,a44790a,a44791a,a44794a,a44797a,a44798a,a44799a,a44802a,a44805a,a44806a,a44809a,a44812a,a44813a,a44814a,a44817a,a44820a,a44821a,a44824a,a44827a,a44828a,a44829a,a44832a,a44835a,a44836a,a44839a,a44842a,a44843a,a44844a,a44847a,a44850a,a44851a,a44854a,a44857a,a44858a,a44859a,a44862a,a44865a,a44866a,a44869a,a44872a,a44873a,a44874a,a44877a,a44880a,a44881a,a44884a,a44887a,a44888a,a44889a,a44892a,a44895a,a44896a,a44899a,a44902a,a44903a,a44904a,a44907a,a44910a,a44911a,a44914a,a44917a,a44918a,a44919a,a44922a,a44925a,a44926a,a44929a,a44932a,a44933a,a44934a,a44937a,a44940a,a44941a,a44944a,a44947a,a44948a,a44949a,a44952a,a44955a,a44956a,a44959a,a44962a,a44963a,a44964a,a44967a,a44970a,a44971a,a44974a,a44977a,a44978a,a44979a,a44982a,a44985a,a44986a,a44989a,a44992a,a44993a,a44994a,a44997a,a45000a,a45001a,a45004a,a45007a,a45008a,a45009a,a45012a,a45015a,a45016a,a45019a,a45022a,a45023a,a45024a,a45027a,a45030a,a45031a,a45034a,a45037a,a45038a,a45039a,a45042a,a45045a,a45046a,a45049a,a45052a,a45053a,a45054a,a45057a,a45060a,a45061a,a45064a,a45067a,a45068a,a45069a,a45072a,a45075a,a45076a,a45079a,a45082a,a45083a,a45084a,a45087a,a45090a,a45091a,a45094a,a45097a,a45098a,a45099a,a45102a,a45105a,a45106a,a45109a,a45112a,a45113a,a45114a,a45117a,a45120a,a45121a,a45124a,a45127a,a45128a,a45129a,a45132a,a45135a,a45136a,a45139a,a45142a,a45143a,a45144a,a45147a,a45150a,a45151a,a45154a,a45157a,a45158a,a45159a,a45162a,a45165a,a45166a,a45169a,a45172a,a45173a,a45174a,a45177a,a45180a,a45181a,a45184a,a45187a,a45188a,a45189a,a45192a,a45195a,a45196a,a45199a,a45202a,a45203a,a45204a,a45207a,a45210a,a45211a,a45214a,a45217a,a45218a,a45219a,a45222a,a45225a,a45226a,a45229a,a45232a,a45233a,a45234a,a45237a,a45240a,a45241a,a45244a,a45247a,a45248a,a45249a,a45252a,a45255a,a45256a,a45259a,a45262a,a45263a,a45264a,a45267a,a45270a,a45271a,a45274a,a45277a,a45278a,a45279a,a45282a,a45285a,a45286a,a45289a,a45292a,a45293a,a45294a,a45297a,a45300a,a45301a,a45304a,a45307a,a45308a,a45309a,a45312a,a45315a,a45316a,a45319a,a45322a,a45323a,a45324a,a45327a,a45330a,a45331a,a45334a,a45337a,a45338a,a45339a,a45342a,a45345a,a45346a,a45349a,a45352a,a45353a,a45354a,a45357a,a45360a,a45361a,a45364a,a45367a,a45368a,a45369a,a45372a,a45375a,a45376a,a45379a,a45382a,a45383a,a45384a,a45387a,a45390a,a45391a,a45394a,a45397a,a45398a,a45399a,a45402a,a45405a,a45406a,a45409a,a45412a,a45413a,a45414a,a45417a,a45420a,a45421a,a45424a,a45427a,a45428a,a45429a,a45432a,a45435a,a45436a,a45439a,a45442a,a45443a,a45444a,a45447a,a45450a,a45451a,a45454a,a45457a,a45458a,a45459a,a45462a,a45465a,a45466a,a45469a,a45472a,a45473a,a45474a,a45477a,a45480a,a45481a,a45484a,a45487a,a45488a,a45489a,a45492a,a45495a,a45496a,a45499a,a45502a,a45503a,a45504a,a45507a,a45510a,a45511a,a45514a,a45517a,a45518a,a45519a,a45522a,a45525a,a45526a,a45529a,a45532a,a45533a,a45534a,a45537a,a45540a,a45541a,a45544a,a45547a,a45548a,a45549a,a45552a,a45555a,a45556a,a45559a,a45562a,a45563a,a45564a,a45567a,a45570a,a45571a,a45574a,a45577a,a45578a,a45579a,a45582a,a45585a,a45586a,a45589a,a45592a,a45593a,a45594a,a45597a,a45600a,a45601a,a45604a,a45607a,a45608a,a45609a,a45612a,a45615a,a45616a,a45619a,a45622a,a45623a,a45624a,a45627a,a45630a,a45631a,a45634a,a45637a,a45638a,a45639a,a45642a,a45645a,a45646a,a45649a,a45652a,a45653a,a45654a,a45657a,a45660a,a45661a,a45664a,a45667a,a45668a,a45669a,a45672a,a45675a,a45676a,a45679a,a45682a,a45683a,a45684a,a45687a,a45690a,a45691a,a45694a,a45697a,a45698a,a45699a,a45702a,a45705a,a45706a,a45709a,a45712a,a45713a,a45714a,a45717a,a45720a,a45721a,a45724a,a45727a,a45728a,a45729a,a45732a,a45735a,a45736a,a45739a,a45742a,a45743a,a45744a,a45747a,a45750a,a45751a,a45754a,a45757a,a45758a,a45759a,a45762a,a45765a,a45766a,a45769a,a45772a,a45773a,a45774a,a45777a,a45780a,a45781a,a45784a,a45787a,a45788a,a45789a,a45792a,a45795a,a45796a,a45799a,a45802a,a45803a,a45804a,a45807a,a45810a,a45811a,a45814a,a45817a,a45818a,a45819a,a45822a,a45825a,a45826a,a45829a,a45832a,a45833a,a45834a,a45837a,a45840a,a45841a,a45844a,a45847a,a45848a,a45849a,a45852a,a45855a,a45856a,a45859a,a45862a,a45863a,a45864a,a45867a,a45870a,a45871a,a45874a,a45877a,a45878a,a45879a,a45882a,a45885a,a45886a,a45889a,a45892a,a45893a,a45894a,a45897a,a45900a,a45901a,a45904a,a45907a,a45908a,a45909a,a45912a,a45915a,a45916a,a45919a,a45922a,a45923a,a45924a,a45927a,a45930a,a45931a,a45934a,a45937a,a45938a,a45939a,a45942a,a45945a,a45946a,a45949a,a45952a,a45953a,a45954a,a45957a,a45960a,a45961a,a45964a,a45967a,a45968a,a45969a,a45972a,a45975a,a45976a,a45979a,a45982a,a45983a,a45984a,a45987a,a45990a,a45991a,a45994a,a45997a,a45998a,a45999a,a46002a,a46005a,a46006a,a46009a,a46012a,a46013a,a46014a,a46017a,a46020a,a46021a,a46024a,a46027a,a46028a,a46029a,a46032a,a46035a,a46036a,a46039a,a46042a,a46043a,a46044a,a46047a,a46050a,a46051a,a46054a,a46057a,a46058a,a46059a,a46062a,a46065a,a46066a,a46069a,a46072a,a46073a,a46074a,a46077a,a46080a,a46081a,a46084a,a46087a,a46088a,a46089a,a46092a,a46095a,a46096a,a46099a,a46102a,a46103a,a46104a,a46107a,a46110a,a46111a,a46114a,a46117a,a46118a,a46119a,a46122a,a46125a,a46126a,a46129a,a46132a,a46133a,a46134a,a46137a,a46140a,a46141a,a46144a,a46147a,a46148a,a46149a,a46152a,a46155a,a46156a,a46159a,a46162a,a46163a,a46164a,a46167a,a46170a,a46171a,a46174a,a46177a,a46178a,a46179a,a46182a,a46185a,a46186a,a46189a,a46192a,a46193a,a46194a,a46197a,a46200a,a46201a,a46204a,a46207a,a46208a,a46209a,a46212a,a46215a,a46216a,a46219a,a46222a,a46223a,a46224a,a46227a,a46230a,a46231a,a46234a,a46237a,a46238a,a46239a,a46242a,a46245a,a46246a,a46249a,a46252a,a46253a,a46254a,a46257a,a46260a,a46261a,a46264a,a46267a,a46268a,a46269a,a46272a,a46275a,a46276a,a46279a,a46282a,a46283a,a46284a,a46287a,a46290a,a46291a,a46294a,a46297a,a46298a,a46299a,a46302a,a46305a,a46306a,a46309a,a46312a,a46313a,a46314a,a46317a,a46320a,a46321a,a46324a,a46327a,a46328a,a46329a,a46332a,a46335a,a46336a,a46339a,a46342a,a46343a,a46344a,a46347a,a46350a,a46351a,a46354a,a46357a,a46358a,a46359a,a46362a,a46365a,a46366a,a46369a,a46372a,a46373a,a46374a,a46377a,a46380a,a46381a,a46384a,a46387a,a46388a,a46389a,a46392a,a46395a,a46396a,a46399a,a46402a,a46403a,a46404a,a46407a,a46410a,a46411a,a46414a,a46417a,a46418a,a46419a,a46422a,a46425a,a46426a,a46429a,a46432a,a46433a,a46434a,a46437a,a46440a,a46441a,a46444a,a46447a,a46448a,a46449a,a46452a,a46455a,a46456a,a46459a,a46462a,a46463a,a46464a,a46467a,a46470a,a46471a,a46474a,a46477a,a46478a,a46479a,a46482a,a46485a,a46486a,a46489a,a46492a,a46493a,a46494a,a46497a,a46500a,a46501a,a46504a,a46507a,a46508a,a46509a,a46512a,a46515a,a46516a,a46519a,a46522a,a46523a,a46524a,a46527a,a46530a,a46531a,a46534a,a46537a,a46538a,a46539a,a46542a,a46545a,a46546a,a46549a,a46552a,a46553a,a46554a,a46557a,a46560a,a46561a,a46564a,a46567a,a46568a,a46569a,a46572a,a46575a,a46576a,a46579a,a46582a,a46583a,a46584a,a46587a,a46590a,a46591a,a46594a,a46597a,a46598a,a46599a,a46602a,a46605a,a46606a,a46609a,a46612a,a46613a,a46614a,a46617a,a46620a,a46621a,a46624a,a46627a,a46628a,a46629a,a46632a,a46635a,a46636a,a46639a,a46642a,a46643a,a46644a,a46647a,a46650a,a46651a,a46654a,a46657a,a46658a,a46659a,a46662a,a46665a,a46666a,a46669a,a46672a,a46673a,a46674a,a46677a,a46680a,a46681a,a46684a,a46687a,a46688a,a46689a,a46692a,a46695a,a46696a,a46699a,a46702a,a46703a,a46704a,a46707a,a46710a,a46711a,a46714a,a46717a,a46718a,a46719a,a46722a,a46725a,a46726a,a46729a,a46732a,a46733a,a46734a,a46737a,a46740a,a46741a,a46744a,a46747a,a46748a,a46749a,a46752a,a46755a,a46756a,a46759a,a46762a,a46763a,a46764a,a46767a,a46770a,a46771a,a46774a,a46777a,a46778a,a46779a,a46782a,a46785a,a46786a,a46789a,a46792a,a46793a,a46794a,a46797a,a46800a,a46801a,a46804a,a46807a,a46808a,a46809a,a46812a,a46815a,a46816a,a46819a,a46822a,a46823a,a46824a,a46827a,a46830a,a46831a,a46834a,a46837a,a46838a,a46839a,a46842a,a46845a,a46846a,a46849a,a46852a,a46853a,a46854a,a46857a,a46860a,a46861a,a46864a,a46867a,a46868a,a46869a,a46872a,a46875a,a46876a,a46879a,a46882a,a46883a,a46884a,a46887a,a46890a,a46891a,a46894a,a46897a,a46898a,a46899a,a46902a,a46905a,a46906a,a46909a,a46912a,a46913a,a46914a,a46917a,a46920a,a46921a,a46924a,a46927a,a46928a,a46929a,a46932a,a46935a,a46936a,a46939a,a46942a,a46943a,a46944a,a46947a,a46950a,a46951a,a46954a,a46957a,a46958a,a46959a,a46962a,a46965a,a46966a,a46969a,a46972a,a46973a,a46974a,a46977a,a46980a,a46981a,a46984a,a46987a,a46988a,a46989a,a46992a,a46995a,a46996a,a46999a,a47002a,a47003a,a47004a,a47007a,a47010a,a47011a,a47014a,a47017a,a47018a,a47019a,a47022a,a47025a,a47026a,a47029a,a47032a,a47033a,a47034a,a47037a,a47040a,a47041a,a47044a,a47047a,a47048a,a47049a,a47052a,a47055a,a47056a,a47059a,a47062a,a47063a,a47064a,a47067a,a47070a,a47071a,a47074a,a47077a,a47078a,a47079a,a47082a,a47085a,a47086a,a47089a,a47092a,a47093a,a47094a,a47097a,a47100a,a47101a,a47104a,a47107a,a47108a,a47109a,a47112a,a47115a,a47116a,a47119a,a47122a,a47123a,a47124a,a47127a,a47130a,a47131a,a47134a,a47137a,a47138a,a47139a,a47142a,a47145a,a47146a,a47149a,a47152a,a47153a,a47154a,a47157a,a47160a,a47161a,a47164a,a47167a,a47168a,a47169a,a47172a,a47175a,a47176a,a47179a,a47182a,a47183a,a47184a,a47187a,a47190a,a47191a,a47194a,a47197a,a47198a,a47199a,a47202a,a47205a,a47206a,a47209a,a47212a,a47213a,a47214a,a47217a,a47220a,a47221a,a47224a,a47227a,a47228a,a47229a,a47232a,a47235a,a47236a,a47239a,a47242a,a47243a,a47244a,a47247a,a47250a,a47251a,a47254a,a47257a,a47258a,a47259a,a47262a,a47265a,a47266a,a47269a,a47272a,a47273a,a47274a,a47277a,a47280a,a47281a,a47284a,a47287a,a47288a,a47289a,a47292a,a47295a,a47296a,a47299a,a47302a,a47303a,a47304a,a47307a,a47310a,a47311a,a47314a,a47317a,a47318a,a47319a,a47322a,a47325a,a47326a,a47329a,a47332a,a47333a,a47334a,a47337a,a47340a,a47341a,a47344a,a47347a,a47348a,a47349a,a47352a,a47355a,a47356a,a47359a,a47362a,a47363a,a47364a,a47367a,a47370a,a47371a,a47374a,a47377a,a47378a,a47379a,a47382a,a47385a,a47386a,a47389a,a47392a,a47393a,a47394a,a47397a,a47400a,a47401a,a47404a,a47407a,a47408a,a47409a,a47412a,a47415a,a47416a,a47419a,a47422a,a47423a,a47424a,a47427a,a47430a,a47431a,a47434a,a47437a,a47438a,a47439a,a47442a,a47445a,a47446a,a47449a,a47452a,a47453a,a47454a,a47457a,a47460a,a47461a,a47464a,a47467a,a47468a,a47469a,a47472a,a47475a,a47476a,a47479a,a47482a,a47483a,a47484a,a47487a,a47490a,a47491a,a47494a,a47497a,a47498a,a47499a,a47502a,a47505a,a47506a,a47509a,a47512a,a47513a,a47514a,a47517a,a47520a,a47521a,a47524a,a47527a,a47528a,a47529a,a47532a,a47535a,a47536a,a47539a,a47542a,a47543a,a47544a,a47547a,a47550a,a47551a,a47554a,a47557a,a47558a,a47559a,a47562a,a47565a,a47566a,a47569a,a47572a,a47573a,a47574a,a47577a,a47580a,a47581a,a47584a,a47587a,a47588a,a47589a,a47592a,a47595a,a47596a,a47599a,a47602a,a47603a,a47604a,a47607a,a47610a,a47611a,a47614a,a47617a,a47618a,a47619a,a47622a,a47625a,a47626a,a47629a,a47632a,a47633a,a47634a,a47637a,a47640a,a47641a,a47644a,a47647a,a47648a,a47649a,a47652a,a47655a,a47656a,a47659a,a47662a,a47663a,a47664a,a47667a,a47670a,a47671a,a47674a,a47677a,a47678a,a47679a,a47682a,a47685a,a47686a,a47689a,a47692a,a47693a,a47694a,a47697a,a47700a,a47701a,a47704a,a47707a,a47708a,a47709a,a47712a,a47715a,a47716a,a47719a,a47722a,a47723a,a47724a,a47727a,a47730a,a47731a,a47734a,a47737a,a47738a,a47739a,a47742a,a47745a,a47746a,a47749a,a47752a,a47753a,a47754a,a47757a,a47760a,a47761a,a47764a,a47767a,a47768a,a47769a,a47772a,a47775a,a47776a,a47779a,a47782a,a47783a,a47784a,a47787a,a47790a,a47791a,a47794a,a47797a,a47798a,a47799a,a47802a,a47805a,a47806a,a47809a,a47812a,a47813a,a47814a,a47817a,a47820a,a47821a,a47824a,a47827a,a47828a,a47829a,a47832a,a47835a,a47836a,a47839a,a47842a,a47843a,a47844a,a47847a,a47850a,a47851a,a47854a,a47857a,a47858a,a47859a,a47862a,a47865a,a47866a,a47869a,a47872a,a47873a,a47874a,a47877a,a47880a,a47881a,a47884a,a47887a,a47888a,a47889a,a47892a,a47895a,a47896a,a47899a,a47902a,a47903a,a47904a,a47907a,a47910a,a47911a,a47914a,a47917a,a47918a,a47919a,a47922a,a47925a,a47926a,a47929a,a47932a,a47933a,a47934a,a47937a,a47940a,a47941a,a47944a,a47947a,a47948a,a47949a,a47952a,a47955a,a47956a,a47959a,a47962a,a47963a,a47964a,a47967a,a47970a,a47971a,a47974a,a47977a,a47978a,a47979a,a47982a,a47985a,a47986a,a47989a,a47992a,a47993a,a47994a,a47997a,a48000a,a48001a,a48004a,a48007a,a48008a,a48009a,a48012a,a48015a,a48016a,a48019a,a48022a,a48023a,a48024a,a48027a,a48030a,a48031a,a48034a,a48037a,a48038a,a48039a,a48042a,a48045a,a48046a,a48049a,a48052a,a48053a,a48054a,a48057a,a48060a,a48061a,a48064a,a48067a,a48068a,a48069a,a48072a,a48075a,a48076a,a48079a,a48082a,a48083a,a48084a,a48087a,a48090a,a48091a,a48094a,a48097a,a48098a,a48099a,a48102a,a48105a,a48106a,a48109a,a48112a,a48113a,a48114a,a48117a,a48120a,a48121a,a48124a,a48127a,a48128a,a48129a,a48132a,a48135a,a48136a,a48139a,a48142a,a48143a,a48144a,a48147a,a48150a,a48151a,a48154a,a48157a,a48158a,a48159a,a48162a,a48165a,a48166a,a48169a,a48172a,a48173a,a48174a,a48177a,a48180a,a48181a,a48184a,a48187a,a48188a,a48189a,a48192a,a48195a,a48196a,a48199a,a48202a,a48203a,a48204a,a48207a,a48210a,a48211a,a48214a,a48217a,a48218a,a48219a,a48222a,a48225a,a48226a,a48229a,a48232a,a48233a,a48234a,a48237a,a48240a,a48241a,a48244a,a48247a,a48248a,a48249a,a48252a,a48255a,a48256a,a48259a,a48262a,a48263a,a48264a,a48267a,a48270a,a48271a,a48274a,a48277a,a48278a,a48279a,a48282a,a48285a,a48286a,a48289a,a48292a,a48293a,a48294a,a48297a,a48300a,a48301a,a48304a,a48307a,a48308a,a48309a,a48312a,a48315a,a48316a,a48319a,a48322a,a48323a,a48324a,a48327a,a48330a,a48331a,a48334a,a48337a,a48338a,a48339a,a48342a,a48345a,a48346a,a48349a,a48352a,a48353a,a48354a,a48357a,a48360a,a48361a,a48364a,a48367a,a48368a,a48369a,a48372a,a48375a,a48376a,a48379a,a48382a,a48383a,a48384a,a48387a,a48390a,a48391a,a48394a,a48397a,a48398a,a48399a,a48402a,a48405a,a48406a,a48409a,a48412a,a48413a,a48414a,a48417a,a48420a,a48421a,a48424a,a48427a,a48428a,a48429a,a48432a,a48435a,a48436a,a48439a,a48442a,a48443a,a48444a,a48447a,a48450a,a48451a,a48454a,a48457a,a48458a,a48459a,a48462a,a48465a,a48466a,a48469a,a48472a,a48473a,a48474a,a48477a,a48480a,a48481a,a48484a,a48487a,a48488a,a48489a,a48492a,a48495a,a48496a,a48499a,a48502a,a48503a,a48504a,a48507a,a48510a,a48511a,a48514a,a48517a,a48518a,a48519a,a48522a,a48525a,a48526a,a48529a,a48532a,a48533a,a48534a,a48537a,a48540a,a48541a,a48544a,a48547a,a48548a,a48549a,a48552a,a48555a,a48556a,a48559a,a48562a,a48563a,a48564a,a48567a,a48570a,a48571a,a48574a,a48577a,a48578a,a48579a,a48582a,a48585a,a48586a,a48589a,a48592a,a48593a,a48594a,a48597a,a48600a,a48601a,a48604a,a48607a,a48608a,a48609a,a48612a,a48615a,a48616a,a48619a,a48622a,a48623a,a48624a,a48627a,a48630a,a48631a,a48634a,a48637a,a48638a,a48639a,a48642a,a48645a,a48646a,a48649a,a48652a,a48653a,a48654a,a48657a,a48660a,a48661a,a48664a,a48667a,a48668a,a48669a,a48672a,a48675a,a48676a,a48679a,a48682a,a48683a,a48684a,a48687a,a48690a,a48691a,a48694a,a48697a,a48698a,a48699a,a48702a,a48705a,a48706a,a48709a,a48712a,a48713a,a48714a,a48717a,a48720a,a48721a,a48724a,a48727a,a48728a,a48729a,a48732a,a48735a,a48736a,a48739a,a48742a,a48743a,a48744a,a48747a,a48750a,a48751a,a48754a,a48757a,a48758a,a48759a,a48762a,a48765a,a48766a,a48769a,a48772a,a48773a,a48774a,a48777a,a48780a,a48781a,a48784a,a48787a,a48788a,a48789a,a48792a,a48795a,a48796a,a48799a,a48802a,a48803a,a48804a,a48807a,a48810a,a48811a,a48814a,a48817a,a48818a,a48819a,a48822a,a48825a,a48826a,a48829a,a48832a,a48833a,a48834a,a48837a,a48840a,a48841a,a48844a,a48847a,a48848a,a48849a,a48852a,a48855a,a48856a,a48859a,a48862a,a48863a,a48864a,a48867a,a48870a,a48871a,a48874a,a48877a,a48878a,a48879a,a48882a,a48885a,a48886a,a48889a,a48892a,a48893a,a48894a,a48897a,a48900a,a48901a,a48904a,a48907a,a48908a,a48909a,a48912a,a48915a,a48916a,a48919a,a48922a,a48923a,a48924a,a48927a,a48930a,a48931a,a48934a,a48937a,a48938a,a48939a,a48942a,a48945a,a48946a,a48949a,a48952a,a48953a,a48954a,a48957a,a48960a,a48961a,a48964a,a48967a,a48968a,a48969a,a48972a,a48975a,a48976a,a48979a,a48982a,a48983a,a48984a,a48987a,a48990a,a48991a,a48994a,a48997a,a48998a,a48999a,a49002a,a49005a,a49006a,a49009a,a49012a,a49013a,a49014a,a49017a,a49020a,a49021a,a49024a,a49027a,a49028a,a49029a,a49032a,a49035a,a49036a,a49039a,a49042a,a49043a,a49044a,a49047a,a49050a,a49051a,a49054a,a49057a,a49058a,a49059a,a49062a,a49065a,a49066a,a49069a,a49072a,a49073a,a49074a,a49077a,a49080a,a49081a,a49084a,a49087a,a49088a,a49089a,a49092a,a49095a,a49096a,a49099a,a49102a,a49103a,a49104a,a49107a,a49110a,a49111a,a49114a,a49117a,a49118a,a49119a,a49122a,a49125a,a49126a,a49129a,a49132a,a49133a,a49134a,a49137a,a49140a,a49141a,a49144a,a49147a,a49148a,a49149a,a49152a,a49155a,a49156a,a49159a,a49162a,a49163a,a49164a,a49167a,a49170a,a49171a,a49174a,a49177a,a49178a,a49179a,a49182a,a49185a,a49186a,a49189a,a49192a,a49193a,a49194a,a49197a,a49200a,a49201a,a49204a,a49207a,a49208a,a49209a,a49212a,a49215a,a49216a,a49219a,a49222a,a49223a,a49224a,a49227a,a49230a,a49231a,a49234a,a49237a,a49238a,a49239a,a49242a,a49245a,a49246a,a49249a,a49252a,a49253a,a49254a,a49257a,a49260a,a49261a,a49264a,a49267a,a49268a,a49269a,a49272a,a49275a,a49276a,a49279a,a49282a,a49283a,a49284a,a49287a,a49290a,a49291a,a49294a,a49297a,a49298a,a49299a,a49302a,a49305a,a49306a,a49309a,a49312a,a49313a,a49314a,a49317a,a49320a,a49321a,a49324a,a49327a,a49328a,a49329a,a49332a,a49335a,a49336a,a49339a,a49342a,a49343a,a49344a,a49347a,a49350a,a49351a,a49354a,a49357a,a49358a,a49359a,a49362a,a49365a,a49366a,a49369a,a49372a,a49373a,a49374a,a49377a,a49380a,a49381a,a49384a,a49387a,a49388a,a49389a,a49392a,a49395a,a49396a,a49399a,a49402a,a49403a,a49404a,a49407a,a49410a,a49411a,a49414a,a49417a,a49418a,a49419a,a49422a,a49425a,a49426a,a49429a,a49432a,a49433a,a49434a,a49437a,a49440a,a49441a,a49444a,a49447a,a49448a,a49449a,a49452a,a49455a,a49456a,a49459a,a49462a,a49463a,a49464a,a49467a,a49470a,a49471a,a49474a,a49477a,a49478a,a49479a,a49482a,a49485a,a49486a,a49489a,a49492a,a49493a,a49494a,a49497a,a49500a,a49501a,a49504a,a49507a,a49508a,a49509a,a49512a,a49515a,a49516a,a49519a,a49522a,a49523a,a49524a,a49527a,a49530a,a49531a,a49534a,a49537a,a49538a,a49539a,a49542a,a49545a,a49546a,a49549a,a49552a,a49553a,a49554a,a49557a,a49560a,a49561a,a49564a,a49567a,a49568a,a49569a,a49572a,a49575a,a49576a,a49579a,a49582a,a49583a,a49584a,a49587a,a49590a,a49591a,a49594a,a49597a,a49598a,a49599a,a49602a,a49605a,a49606a,a49609a,a49612a,a49613a,a49614a,a49617a,a49620a,a49621a,a49624a,a49627a,a49628a,a49629a,a49632a,a49635a,a49636a,a49639a,a49642a,a49643a,a49644a,a49647a,a49650a,a49651a,a49654a,a49657a,a49658a,a49659a,a49662a,a49665a,a49666a,a49669a,a49672a,a49673a,a49674a,a49677a,a49680a,a49681a,a49684a,a49687a,a49688a,a49689a,a49692a,a49695a,a49696a,a49699a,a49702a,a49703a,a49704a,a49707a,a49710a,a49711a,a49714a,a49717a,a49718a,a49719a,a49722a,a49725a,a49726a,a49729a,a49732a,a49733a,a49734a,a49737a,a49740a,a49741a,a49744a,a49747a,a49748a,a49749a,a49752a,a49755a,a49756a,a49759a,a49762a,a49763a,a49764a,a49767a,a49770a,a49771a,a49774a,a49777a,a49778a,a49779a,a49782a,a49785a,a49786a,a49789a,a49792a,a49793a,a49794a,a49797a,a49800a,a49801a,a49804a,a49807a,a49808a,a49809a,a49812a,a49815a,a49816a,a49819a,a49822a,a49823a,a49824a,a49827a,a49830a,a49831a,a49834a,a49837a,a49838a,a49839a,a49842a,a49845a,a49846a,a49849a,a49852a,a49853a,a49854a,a49857a,a49860a,a49861a,a49864a,a49867a,a49868a,a49869a,a49872a,a49875a,a49876a,a49879a,a49882a,a49883a,a49884a,a49887a,a49890a,a49891a,a49894a,a49897a,a49898a,a49899a,a49902a,a49905a,a49906a,a49909a,a49912a,a49913a,a49914a,a49917a,a49920a,a49921a,a49924a,a49927a,a49928a,a49929a,a49932a,a49935a,a49936a,a49939a,a49942a,a49943a,a49944a,a49947a,a49950a,a49951a,a49954a,a49957a,a49958a,a49959a,a49962a,a49965a,a49966a,a49969a,a49972a,a49973a,a49974a,a49977a,a49980a,a49981a,a49984a,a49987a,a49988a,a49989a,a49992a,a49995a,a49996a,a49999a,a50002a,a50003a,a50004a,a50007a,a50010a,a50011a,a50014a,a50017a,a50018a,a50019a,a50022a,a50025a,a50026a,a50029a,a50032a,a50033a,a50034a,a50037a,a50040a,a50041a,a50044a,a50047a,a50048a,a50049a,a50052a,a50055a,a50056a,a50059a,a50062a,a50063a,a50064a,a50067a,a50070a,a50071a,a50074a,a50077a,a50078a,a50079a,a50082a,a50085a,a50086a,a50089a,a50092a,a50093a,a50094a,a50097a,a50100a,a50101a,a50104a,a50107a,a50108a,a50109a,a50112a,a50115a,a50116a,a50119a,a50122a,a50123a,a50124a,a50127a,a50130a,a50131a,a50134a,a50137a,a50138a,a50139a,a50142a,a50145a,a50146a,a50149a,a50152a,a50153a,a50154a,a50157a,a50160a,a50161a,a50164a,a50167a,a50168a,a50169a,a50172a,a50175a,a50176a,a50179a,a50182a,a50183a,a50184a,a50187a,a50190a,a50191a,a50194a,a50197a,a50198a,a50199a,a50202a,a50205a,a50206a,a50209a,a50212a,a50213a,a50214a,a50217a,a50220a,a50221a,a50224a,a50227a,a50228a,a50229a,a50232a,a50235a,a50236a,a50239a,a50242a,a50243a,a50244a,a50247a,a50250a,a50251a,a50254a,a50257a,a50258a,a50259a,a50262a,a50265a,a50266a,a50269a,a50272a,a50273a,a50274a,a50277a,a50280a,a50281a,a50284a,a50287a,a50288a,a50289a,a50292a,a50295a,a50296a,a50299a,a50302a,a50303a,a50304a,a50307a,a50310a,a50311a,a50314a,a50317a,a50318a,a50319a,a50322a,a50325a,a50326a,a50329a,a50332a,a50333a,a50334a,a50337a,a50340a,a50341a,a50344a,a50347a,a50348a,a50349a,a50352a,a50355a,a50356a,a50359a,a50362a,a50363a,a50364a,a50367a,a50370a,a50371a,a50374a,a50377a,a50378a,a50379a,a50382a,a50385a,a50386a,a50389a,a50392a,a50393a,a50394a,a50397a,a50400a,a50401a,a50404a,a50407a,a50408a,a50409a,a50412a,a50415a,a50416a,a50419a,a50422a,a50423a,a50424a,a50427a,a50430a,a50431a,a50434a,a50437a,a50438a,a50439a,a50442a,a50445a,a50446a,a50449a,a50452a,a50453a,a50454a,a50457a,a50460a,a50461a,a50464a,a50467a,a50468a,a50469a,a50472a,a50475a,a50476a,a50479a,a50482a,a50483a,a50484a,a50487a,a50490a,a50491a,a50494a,a50497a,a50498a,a50499a,a50502a,a50505a,a50506a,a50509a,a50512a,a50513a,a50514a,a50517a,a50520a,a50521a,a50524a,a50527a,a50528a,a50529a,a50532a,a50535a,a50536a,a50539a,a50542a,a50543a,a50544a,a50547a,a50550a,a50551a,a50554a,a50557a,a50558a,a50559a,a50562a,a50565a,a50566a,a50569a,a50572a,a50573a,a50574a,a50577a,a50580a,a50581a,a50584a,a50587a,a50588a,a50589a,a50592a,a50595a,a50596a,a50599a,a50602a,a50603a,a50604a,a50607a,a50610a,a50611a,a50614a,a50617a,a50618a,a50619a,a50622a,a50625a,a50626a,a50629a,a50632a,a50633a,a50634a,a50637a,a50640a,a50641a,a50644a,a50647a,a50648a,a50649a,a50652a,a50655a,a50656a,a50659a,a50662a,a50663a,a50664a,a50667a,a50670a,a50671a,a50674a,a50677a,a50678a,a50679a,a50682a,a50685a,a50686a,a50689a,a50692a,a50693a,a50694a,a50697a,a50700a,a50701a,a50704a,a50707a,a50708a,a50709a,a50712a,a50715a,a50716a,a50719a,a50722a,a50723a,a50724a,a50727a,a50730a,a50731a,a50734a,a50737a,a50738a,a50739a,a50742a,a50745a,a50746a,a50749a,a50752a,a50753a,a50754a,a50757a,a50760a,a50761a,a50764a,a50767a,a50768a,a50769a,a50772a,a50775a,a50776a,a50779a,a50782a,a50783a,a50784a,a50787a,a50790a,a50791a,a50794a,a50797a,a50798a,a50799a,a50802a,a50805a,a50806a,a50809a,a50812a,a50813a,a50814a,a50817a,a50820a,a50821a,a50824a,a50827a,a50828a,a50829a,a50832a,a50835a,a50836a,a50839a,a50842a,a50843a,a50844a,a50847a,a50850a,a50851a,a50854a,a50857a,a50858a,a50859a,a50862a,a50865a,a50866a,a50869a,a50872a,a50873a,a50874a,a50877a,a50880a,a50881a,a50884a,a50887a,a50888a,a50889a,a50892a,a50895a,a50896a,a50899a,a50902a,a50903a,a50904a,a50907a,a50910a,a50911a,a50914a,a50917a,a50918a,a50919a,a50922a,a50925a,a50926a,a50929a,a50932a,a50933a,a50934a,a50937a,a50940a,a50941a,a50944a,a50947a,a50948a,a50949a,a50952a,a50955a,a50956a,a50959a,a50962a,a50963a,a50964a,a50967a,a50970a,a50971a,a50974a,a50977a,a50978a,a50979a,a50982a,a50985a,a50986a,a50989a,a50992a,a50993a,a50994a,a50997a,a51000a,a51001a,a51004a,a51007a,a51008a,a51009a,a51012a,a51015a,a51016a,a51019a,a51022a,a51023a,a51024a,a51027a,a51030a,a51031a,a51034a,a51037a,a51038a,a51039a,a51042a,a51045a,a51046a,a51049a,a51052a,a51053a,a51054a,a51057a,a51060a,a51061a,a51064a,a51067a,a51068a,a51069a,a51072a,a51075a,a51076a,a51079a,a51082a,a51083a,a51084a,a51087a,a51090a,a51091a,a51094a,a51097a,a51098a,a51099a,a51102a,a51105a,a51106a,a51109a,a51112a,a51113a,a51114a,a51117a,a51120a,a51121a,a51124a,a51127a,a51128a,a51129a,a51132a,a51135a,a51136a,a51139a,a51142a,a51143a,a51144a,a51147a,a51150a,a51151a,a51154a,a51157a,a51158a,a51159a,a51162a,a51165a,a51166a,a51169a,a51172a,a51173a,a51174a,a51177a,a51180a,a51181a,a51184a,a51187a,a51188a,a51189a,a51192a,a51195a,a51196a,a51199a,a51202a,a51203a,a51204a,a51207a,a51210a,a51211a,a51214a,a51217a,a51218a,a51219a,a51222a,a51225a,a51226a,a51229a,a51232a,a51233a,a51234a,a51237a,a51240a,a51241a,a51244a,a51247a,a51248a,a51249a,a51252a,a51255a,a51256a,a51259a,a51262a,a51263a,a51264a,a51267a,a51270a,a51271a,a51274a,a51277a,a51278a,a51279a,a51282a,a51285a,a51286a,a51289a,a51292a,a51293a,a51294a,a51297a,a51300a,a51301a,a51304a,a51307a,a51308a,a51309a,a51312a,a51315a,a51316a,a51319a,a51322a,a51323a,a51324a,a51327a,a51330a,a51331a,a51334a,a51337a,a51338a,a51339a,a51342a,a51345a,a51346a,a51349a,a51352a,a51353a,a51354a,a51357a,a51360a,a51361a,a51364a,a51367a,a51368a,a51369a,a51372a,a51375a,a51376a,a51379a,a51382a,a51383a,a51384a,a51387a,a51390a,a51391a,a51394a,a51397a,a51398a,a51399a,a51402a,a51405a,a51406a,a51409a,a51412a,a51413a,a51414a,a51417a,a51420a,a51421a,a51424a,a51427a,a51428a,a51429a,a51432a,a51435a,a51436a,a51439a,a51442a,a51443a,a51444a,a51447a,a51450a,a51451a,a51454a,a51457a,a51458a,a51459a,a51462a,a51465a,a51466a,a51469a,a51472a,a51473a,a51474a,a51477a,a51480a,a51481a,a51484a,a51487a,a51488a,a51489a,a51492a,a51495a,a51496a,a51499a,a51502a,a51503a,a51504a,a51507a,a51510a,a51511a,a51514a,a51517a,a51518a,a51519a,a51522a,a51525a,a51526a,a51529a,a51532a,a51533a,a51534a,a51537a,a51540a,a51541a,a51544a,a51547a,a51548a,a51549a,a51552a,a51555a,a51556a,a51559a,a51562a,a51563a,a51564a,a51567a,a51570a,a51571a,a51574a,a51577a,a51578a,a51579a,a51582a,a51585a,a51586a,a51589a,a51592a,a51593a,a51594a,a51597a,a51600a,a51601a,a51604a,a51607a,a51608a,a51609a,a51612a,a51615a,a51616a,a51619a,a51622a,a51623a,a51624a,a51627a,a51630a,a51631a,a51634a,a51637a,a51638a,a51639a,a51642a,a51645a,a51646a,a51649a,a51652a,a51653a,a51654a,a51657a,a51660a,a51661a,a51664a,a51667a,a51668a,a51669a,a51672a,a51675a,a51676a,a51679a,a51682a,a51683a,a51684a,a51687a,a51690a,a51691a,a51694a,a51697a,a51698a,a51699a,a51702a,a51705a,a51706a,a51709a,a51712a,a51713a,a51714a,a51717a,a51720a,a51721a,a51724a,a51727a,a51728a,a51729a,a51732a,a51735a,a51736a,a51739a,a51742a,a51743a,a51744a,a51747a,a51750a,a51751a,a51754a,a51757a,a51758a,a51759a,a51762a,a51765a,a51766a,a51769a,a51773a,a51774a,a51775a,a51776a,a51779a,a51782a,a51783a,a51786a,a51789a,a51790a,a51791a,a51794a,a51797a,a51798a,a51801a,a51805a,a51806a,a51807a,a51808a,a51811a,a51814a,a51815a,a51818a,a51821a,a51822a,a51823a,a51826a,a51829a,a51830a,a51833a,a51837a,a51838a,a51839a,a51840a,a51843a,a51846a,a51847a,a51850a,a51853a,a51854a,a51855a,a51858a,a51861a,a51862a,a51865a,a51869a,a51870a,a51871a,a51872a,a51875a,a51878a,a51879a,a51882a,a51885a,a51886a,a51887a,a51890a,a51893a,a51894a,a51897a,a51901a,a51902a,a51903a,a51904a,a51907a,a51910a,a51911a,a51914a,a51917a,a51918a,a51919a,a51922a,a51925a,a51926a,a51929a,a51933a,a51934a,a51935a,a51936a,a51939a,a51942a,a51943a,a51946a,a51949a,a51950a,a51951a,a51954a,a51957a,a51958a,a51961a,a51965a,a51966a,a51967a,a51968a,a51971a,a51974a,a51975a,a51978a,a51981a,a51982a,a51983a,a51986a,a51989a,a51990a,a51993a,a51997a,a51998a,a51999a,a52000a,a52003a,a52006a,a52007a,a52010a,a52013a,a52014a,a52015a,a52018a,a52021a,a52022a,a52025a,a52029a,a52030a,a52031a,a52032a,a52035a,a52038a,a52039a,a52042a,a52045a,a52046a,a52047a,a52050a,a52053a,a52054a,a52057a,a52061a,a52062a,a52063a,a52064a,a52067a,a52070a,a52071a,a52074a,a52077a,a52078a,a52079a,a52082a,a52085a,a52086a,a52089a,a52093a,a52094a,a52095a,a52096a,a52099a,a52102a,a52103a,a52106a,a52109a,a52110a,a52111a,a52114a,a52117a,a52118a,a52121a,a52125a,a52126a,a52127a,a52128a,a52131a,a52134a,a52135a,a52138a,a52141a,a52142a,a52143a,a52146a,a52149a,a52150a,a52153a,a52157a,a52158a,a52159a,a52160a,a52163a,a52166a,a52167a,a52170a,a52173a,a52174a,a52175a,a52178a,a52181a,a52182a,a52185a,a52189a,a52190a,a52191a,a52192a,a52195a,a52198a,a52199a,a52202a,a52205a,a52206a,a52207a,a52210a,a52213a,a52214a,a52217a,a52221a,a52222a,a52223a,a52224a,a52227a,a52230a,a52231a,a52234a,a52237a,a52238a,a52239a,a52242a,a52245a,a52246a,a52249a,a52253a,a52254a,a52255a,a52256a,a52259a,a52262a,a52263a,a52266a,a52269a,a52270a,a52271a,a52274a,a52277a,a52278a,a52281a,a52285a,a52286a,a52287a,a52288a,a52291a,a52294a,a52295a,a52298a,a52301a,a52302a,a52303a,a52306a,a52309a,a52310a,a52313a,a52317a,a52318a,a52319a,a52320a,a52323a,a52326a,a52327a,a52330a,a52333a,a52334a,a52335a,a52338a,a52341a,a52342a,a52345a,a52349a,a52350a,a52351a,a52352a,a52355a,a52358a,a52359a,a52362a,a52365a,a52366a,a52367a,a52370a,a52373a,a52374a,a52377a,a52381a,a52382a,a52383a,a52384a,a52387a,a52390a,a52391a,a52394a,a52397a,a52398a,a52399a,a52402a,a52405a,a52406a,a52409a,a52413a,a52414a,a52415a,a52416a,a52419a,a52422a,a52423a,a52426a,a52429a,a52430a,a52431a,a52434a,a52437a,a52438a,a52441a,a52445a,a52446a,a52447a,a52448a,a52451a,a52454a,a52455a,a52458a,a52461a,a52462a,a52463a,a52466a,a52469a,a52470a,a52473a,a52477a,a52478a,a52479a,a52480a,a52483a,a52486a,a52487a,a52490a,a52493a,a52494a,a52495a,a52498a,a52501a,a52502a,a52505a,a52509a,a52510a,a52511a,a52512a,a52515a,a52518a,a52519a,a52522a,a52525a,a52526a,a52527a,a52530a,a52533a,a52534a,a52537a,a52541a,a52542a,a52543a,a52544a,a52547a,a52550a,a52551a,a52554a,a52557a,a52558a,a52559a,a52562a,a52565a,a52566a,a52569a,a52573a,a52574a,a52575a,a52576a,a52579a,a52582a,a52583a,a52586a,a52589a,a52590a,a52591a,a52594a,a52597a,a52598a,a52601a,a52605a,a52606a,a52607a,a52608a,a52611a,a52614a,a52615a,a52618a,a52621a,a52622a,a52623a,a52626a,a52629a,a52630a,a52633a,a52637a,a52638a,a52639a,a52640a,a52643a,a52646a,a52647a,a52650a,a52653a,a52654a,a52655a,a52658a,a52661a,a52662a,a52665a,a52669a,a52670a,a52671a,a52672a,a52675a,a52678a,a52679a,a52682a,a52685a,a52686a,a52687a,a52690a,a52693a,a52694a,a52697a,a52701a,a52702a,a52703a,a52704a,a52707a,a52710a,a52711a,a52714a,a52717a,a52718a,a52719a,a52722a,a52725a,a52726a,a52729a,a52733a,a52734a,a52735a,a52736a,a52739a,a52742a,a52743a,a52746a,a52749a,a52750a,a52751a,a52754a,a52757a,a52758a,a52761a,a52765a,a52766a,a52767a,a52768a,a52771a,a52774a,a52775a,a52778a,a52781a,a52782a,a52783a,a52786a,a52789a,a52790a,a52793a,a52797a,a52798a,a52799a,a52800a,a52803a,a52806a,a52807a,a52810a,a52813a,a52814a,a52815a,a52818a,a52821a,a52822a,a52825a,a52829a,a52830a,a52831a,a52832a,a52835a,a52838a,a52839a,a52842a,a52845a,a52846a,a52847a,a52850a,a52853a,a52854a,a52857a,a52861a,a52862a,a52863a,a52864a,a52867a,a52870a,a52871a,a52874a,a52877a,a52878a,a52879a,a52882a,a52885a,a52886a,a52889a,a52893a,a52894a,a52895a,a52896a,a52899a,a52902a,a52903a,a52906a,a52909a,a52910a,a52911a,a52914a,a52917a,a52918a,a52921a,a52925a,a52926a,a52927a,a52928a,a52931a,a52934a,a52935a,a52938a,a52941a,a52942a,a52943a,a52946a,a52949a,a52950a,a52953a,a52957a,a52958a,a52959a,a52960a,a52963a,a52966a,a52967a,a52970a,a52973a,a52974a,a52975a,a52978a,a52981a,a52982a,a52985a,a52989a,a52990a,a52991a,a52992a,a52995a,a52998a,a52999a,a53002a,a53005a,a53006a,a53007a,a53010a,a53013a,a53014a,a53017a,a53021a,a53022a,a53023a,a53024a,a53027a,a53030a,a53031a,a53034a,a53037a,a53038a,a53039a,a53042a,a53045a,a53046a,a53049a,a53053a,a53054a,a53055a,a53056a,a53059a,a53062a,a53063a,a53066a,a53069a,a53070a,a53071a,a53074a,a53077a,a53078a,a53081a,a53085a,a53086a,a53087a,a53088a,a53091a,a53094a,a53095a,a53098a,a53101a,a53102a,a53103a,a53106a,a53109a,a53110a,a53113a,a53117a,a53118a,a53119a,a53120a,a53123a,a53126a,a53127a,a53130a,a53133a,a53134a,a53135a,a53138a,a53141a,a53142a,a53145a,a53149a,a53150a,a53151a,a53152a,a53155a,a53158a,a53159a,a53162a,a53165a,a53166a,a53167a,a53170a,a53173a,a53174a,a53177a,a53181a,a53182a,a53183a,a53184a,a53187a,a53190a,a53191a,a53194a,a53197a,a53198a,a53199a,a53202a,a53205a,a53206a,a53209a,a53213a,a53214a,a53215a,a53216a,a53219a,a53222a,a53223a,a53226a,a53229a,a53230a,a53231a,a53234a,a53237a,a53238a,a53241a,a53245a,a53246a,a53247a,a53248a,a53251a,a53254a,a53255a,a53258a,a53261a,a53262a,a53263a,a53266a,a53269a,a53270a,a53273a,a53277a,a53278a,a53279a,a53280a,a53283a,a53286a,a53287a,a53290a,a53293a,a53294a,a53295a,a53298a,a53301a,a53302a,a53305a,a53309a,a53310a,a53311a,a53312a,a53315a,a53318a,a53319a,a53322a,a53325a,a53326a,a53327a,a53330a,a53333a,a53334a,a53337a,a53341a,a53342a,a53343a,a53344a,a53347a,a53350a,a53351a,a53354a,a53357a,a53358a,a53359a,a53362a,a53365a,a53366a,a53369a,a53373a,a53374a,a53375a,a53376a,a53379a,a53382a,a53383a,a53386a,a53389a,a53390a,a53391a,a53394a,a53397a,a53398a,a53401a,a53405a,a53406a,a53407a,a53408a,a53411a,a53414a,a53415a,a53418a,a53421a,a53422a,a53423a,a53426a,a53429a,a53430a,a53433a,a53437a,a53438a,a53439a,a53440a,a53443a,a53446a,a53447a,a53450a,a53453a,a53454a,a53455a,a53458a,a53461a,a53462a,a53465a,a53469a,a53470a,a53471a,a53472a,a53475a,a53478a,a53479a,a53482a,a53485a,a53486a,a53487a,a53490a,a53493a,a53494a,a53497a,a53501a,a53502a,a53503a,a53504a,a53507a,a53510a,a53511a,a53514a,a53517a,a53518a,a53519a,a53522a,a53525a,a53526a,a53529a,a53533a,a53534a,a53535a,a53536a,a53539a,a53542a,a53543a,a53546a,a53549a,a53550a,a53551a,a53554a,a53557a,a53558a,a53561a,a53565a,a53566a,a53567a,a53568a,a53571a,a53574a,a53575a,a53578a,a53581a,a53582a,a53583a,a53586a,a53589a,a53590a,a53593a,a53597a,a53598a,a53599a,a53600a,a53603a,a53606a,a53607a,a53610a,a53613a,a53614a,a53615a,a53618a,a53621a,a53622a,a53625a,a53629a,a53630a,a53631a,a53632a,a53635a,a53638a,a53639a,a53642a,a53645a,a53646a,a53647a,a53650a,a53653a,a53654a,a53657a,a53661a,a53662a,a53663a,a53664a,a53667a,a53670a,a53671a,a53674a,a53677a,a53678a,a53679a,a53682a,a53685a,a53686a,a53689a,a53693a,a53694a,a53695a,a53696a,a53699a,a53702a,a53703a,a53706a,a53709a,a53710a,a53711a,a53714a,a53717a,a53718a,a53721a,a53725a,a53726a,a53727a,a53728a,a53731a,a53734a,a53735a,a53738a,a53741a,a53742a,a53743a,a53746a,a53749a,a53750a,a53753a,a53757a,a53758a,a53759a,a53760a,a53763a,a53766a,a53767a,a53770a,a53773a,a53774a,a53775a,a53778a,a53781a,a53782a,a53785a,a53789a,a53790a,a53791a,a53792a,a53795a,a53798a,a53799a,a53802a,a53805a,a53806a,a53807a,a53810a,a53813a,a53814a,a53817a,a53821a,a53822a,a53823a,a53824a,a53827a,a53830a,a53831a,a53834a,a53837a,a53838a,a53839a,a53842a,a53845a,a53846a,a53849a,a53853a,a53854a,a53855a,a53856a,a53859a,a53862a,a53863a,a53866a,a53869a,a53870a,a53871a,a53874a,a53877a,a53878a,a53881a,a53885a,a53886a,a53887a,a53888a,a53891a,a53894a,a53895a,a53898a,a53901a,a53902a,a53903a,a53906a,a53909a,a53910a,a53913a,a53917a,a53918a,a53919a,a53920a,a53923a,a53926a,a53927a,a53930a,a53933a,a53934a,a53935a,a53938a,a53941a,a53942a,a53945a,a53949a,a53950a,a53951a,a53952a,a53955a,a53958a,a53959a,a53962a,a53965a,a53966a,a53967a,a53970a,a53973a,a53974a,a53977a,a53981a,a53982a,a53983a,a53984a,a53987a,a53990a,a53991a,a53994a,a53997a,a53998a,a53999a,a54002a,a54005a,a54006a,a54009a,a54013a,a54014a,a54015a,a54016a,a54019a,a54022a,a54023a,a54026a,a54029a,a54030a,a54031a,a54034a,a54037a,a54038a,a54041a,a54045a,a54046a,a54047a,a54048a,a54051a,a54054a,a54055a,a54058a,a54061a,a54062a,a54063a,a54066a,a54069a,a54070a,a54073a,a54077a,a54078a,a54079a,a54080a,a54083a,a54086a,a54087a,a54090a,a54093a,a54094a,a54095a,a54098a,a54101a,a54102a,a54105a,a54109a,a54110a,a54111a,a54112a,a54115a,a54118a,a54119a,a54122a,a54125a,a54126a,a54127a,a54130a,a54133a,a54134a,a54137a,a54141a,a54142a,a54143a,a54144a,a54147a,a54150a,a54151a,a54154a,a54157a,a54158a,a54159a,a54162a,a54165a,a54166a,a54169a,a54173a,a54174a,a54175a,a54176a,a54179a,a54182a,a54183a,a54186a,a54189a,a54190a,a54191a,a54194a,a54197a,a54198a,a54201a,a54205a,a54206a,a54207a,a54208a,a54211a,a54214a,a54215a,a54218a,a54221a,a54222a,a54223a,a54226a,a54229a,a54230a,a54233a,a54237a,a54238a,a54239a,a54240a,a54243a,a54246a,a54247a,a54250a,a54253a,a54254a,a54255a,a54258a,a54261a,a54262a,a54265a,a54269a,a54270a,a54271a,a54272a,a54275a,a54278a,a54279a,a54282a,a54285a,a54286a,a54287a,a54290a,a54293a,a54294a,a54297a,a54301a,a54302a,a54303a,a54304a,a54307a,a54310a,a54311a,a54314a,a54317a,a54318a,a54319a,a54322a,a54325a,a54326a,a54329a,a54333a,a54334a,a54335a,a54336a,a54339a,a54342a,a54343a,a54346a,a54349a,a54350a,a54351a,a54354a,a54357a,a54358a,a54361a,a54365a,a54366a,a54367a,a54368a,a54371a,a54374a,a54375a,a54378a,a54381a,a54382a,a54383a,a54386a,a54389a,a54390a,a54393a,a54397a,a54398a,a54399a,a54400a,a54403a,a54406a,a54407a,a54410a,a54413a,a54414a,a54415a,a54418a,a54421a,a54422a,a54425a,a54429a,a54430a,a54431a,a54432a,a54435a,a54438a,a54439a,a54442a,a54445a,a54446a,a54447a,a54450a,a54453a,a54454a,a54457a,a54461a,a54462a,a54463a,a54464a,a54467a,a54470a,a54471a,a54474a,a54477a,a54478a,a54479a,a54482a,a54485a,a54486a,a54489a,a54493a,a54494a,a54495a,a54496a,a54499a,a54502a,a54503a,a54506a,a54509a,a54510a,a54511a,a54514a,a54517a,a54518a,a54521a,a54525a,a54526a,a54527a,a54528a,a54531a,a54534a,a54535a,a54538a,a54541a,a54542a,a54543a,a54546a,a54549a,a54550a,a54553a,a54557a,a54558a,a54559a,a54560a,a54563a,a54566a,a54567a,a54570a,a54573a,a54574a,a54575a,a54578a,a54581a,a54582a,a54585a,a54589a,a54590a,a54591a,a54592a,a54595a,a54598a,a54599a,a54602a,a54605a,a54606a,a54607a,a54610a,a54613a,a54614a,a54617a,a54621a,a54622a,a54623a,a54624a,a54627a,a54630a,a54631a,a54634a,a54637a,a54638a,a54639a,a54642a,a54645a,a54646a,a54649a,a54653a,a54654a,a54655a,a54656a,a54659a,a54662a,a54663a,a54666a,a54669a,a54670a,a54671a,a54674a,a54677a,a54678a,a54681a,a54685a,a54686a,a54687a,a54688a,a54691a,a54694a,a54695a,a54698a,a54701a,a54702a,a54703a,a54706a,a54709a,a54710a,a54713a,a54717a,a54718a,a54719a,a54720a,a54723a,a54726a,a54727a,a54730a,a54733a,a54734a,a54735a,a54738a,a54741a,a54742a,a54745a,a54749a,a54750a,a54751a,a54752a,a54755a,a54758a,a54759a,a54762a,a54765a,a54766a,a54767a,a54770a,a54773a,a54774a,a54777a,a54781a,a54782a,a54783a,a54784a,a54787a,a54790a,a54791a,a54794a,a54797a,a54798a,a54799a,a54802a,a54805a,a54806a,a54809a,a54813a,a54814a,a54815a,a54816a,a54819a,a54822a,a54823a,a54826a,a54829a,a54830a,a54831a,a54834a,a54837a,a54838a,a54841a,a54845a,a54846a,a54847a,a54848a,a54851a,a54854a,a54855a,a54858a,a54861a,a54862a,a54863a,a54866a,a54869a,a54870a,a54873a,a54877a,a54878a,a54879a,a54880a,a54883a,a54886a,a54887a,a54890a,a54893a,a54894a,a54895a,a54898a,a54901a,a54902a,a54905a,a54909a,a54910a,a54911a,a54912a,a54915a,a54918a,a54919a,a54922a,a54925a,a54926a,a54927a,a54930a,a54933a,a54934a,a54937a,a54941a,a54942a,a54943a,a54944a,a54947a,a54950a,a54951a,a54954a,a54957a,a54958a,a54959a,a54962a,a54965a,a54966a,a54969a,a54973a,a54974a,a54975a,a54976a,a54979a,a54982a,a54983a,a54986a,a54989a,a54990a,a54991a,a54994a,a54997a,a54998a,a55001a,a55005a,a55006a,a55007a,a55008a,a55011a,a55014a,a55015a,a55018a,a55021a,a55022a,a55023a,a55026a,a55029a,a55030a,a55033a,a55037a,a55038a,a55039a,a55040a,a55043a,a55046a,a55047a,a55050a,a55053a,a55054a,a55055a,a55058a,a55061a,a55062a,a55065a,a55069a,a55070a,a55071a,a55072a,a55075a,a55078a,a55079a,a55082a,a55085a,a55086a,a55087a,a55090a,a55093a,a55094a,a55097a,a55101a,a55102a,a55103a,a55104a,a55107a,a55110a,a55111a,a55114a,a55117a,a55118a,a55119a,a55122a,a55125a,a55126a,a55129a,a55133a,a55134a,a55135a,a55136a,a55139a,a55142a,a55143a,a55146a,a55149a,a55150a,a55151a,a55154a,a55157a,a55158a,a55161a,a55165a,a55166a,a55167a,a55168a,a55171a,a55174a,a55175a,a55178a,a55181a,a55182a,a55183a,a55186a,a55189a,a55190a,a55193a,a55197a,a55198a,a55199a,a55200a,a55203a,a55206a,a55207a,a55210a,a55213a,a55214a,a55215a,a55218a,a55221a,a55222a,a55225a,a55229a,a55230a,a55231a,a55232a,a55235a,a55238a,a55239a,a55242a,a55245a,a55246a,a55247a,a55250a,a55253a,a55254a,a55257a,a55261a,a55262a,a55263a,a55264a,a55267a,a55270a,a55271a,a55274a,a55277a,a55278a,a55279a,a55282a,a55285a,a55286a,a55289a,a55293a,a55294a,a55295a,a55296a,a55299a,a55302a,a55303a,a55306a,a55309a,a55310a,a55311a,a55314a,a55317a,a55318a,a55321a,a55325a,a55326a,a55327a,a55328a,a55331a,a55334a,a55335a,a55338a,a55341a,a55342a,a55343a,a55346a,a55349a,a55350a,a55353a,a55357a,a55358a,a55359a,a55360a,a55363a,a55366a,a55367a,a55370a,a55373a,a55374a,a55375a,a55378a,a55381a,a55382a,a55385a,a55389a,a55390a,a55391a,a55392a,a55395a,a55398a,a55399a,a55402a,a55405a,a55406a,a55407a,a55410a,a55413a,a55414a,a55417a,a55421a,a55422a,a55423a,a55424a,a55427a,a55430a,a55431a,a55434a,a55437a,a55438a,a55439a,a55442a,a55445a,a55446a,a55449a,a55453a,a55454a,a55455a,a55456a,a55459a,a55462a,a55463a,a55466a,a55469a,a55470a,a55471a,a55474a,a55477a,a55478a,a55481a,a55485a,a55486a,a55487a,a55488a,a55491a,a55494a,a55495a,a55498a,a55501a,a55502a,a55503a,a55506a,a55509a,a55510a,a55513a,a55517a,a55518a,a55519a,a55520a,a55523a,a55526a,a55527a,a55530a,a55533a,a55534a,a55535a,a55538a,a55541a,a55542a,a55545a,a55549a,a55550a,a55551a,a55552a,a55555a,a55558a,a55559a,a55562a,a55565a,a55566a,a55567a,a55570a,a55573a,a55574a,a55577a,a55581a,a55582a,a55583a,a55584a,a55587a,a55590a,a55591a,a55594a,a55597a,a55598a,a55599a,a55602a,a55605a,a55606a,a55609a,a55613a,a55614a,a55615a,a55616a,a55619a,a55622a,a55623a,a55626a,a55629a,a55630a,a55631a,a55634a,a55637a,a55638a,a55641a,a55645a,a55646a,a55647a,a55648a,a55651a,a55654a,a55655a,a55658a,a55661a,a55662a,a55663a,a55666a,a55669a,a55670a,a55673a,a55677a,a55678a,a55679a,a55680a,a55683a,a55686a,a55687a,a55690a,a55693a,a55694a,a55695a,a55698a,a55701a,a55702a,a55705a,a55709a,a55710a,a55711a,a55712a,a55715a,a55718a,a55719a,a55722a,a55725a,a55726a,a55727a,a55730a,a55733a,a55734a,a55737a,a55741a,a55742a,a55743a,a55744a,a55747a,a55750a,a55751a,a55754a,a55757a,a55758a,a55759a,a55762a,a55765a,a55766a,a55769a,a55773a,a55774a,a55775a,a55776a,a55779a,a55782a,a55783a,a55786a,a55789a,a55790a,a55791a,a55794a,a55797a,a55798a,a55801a,a55805a,a55806a,a55807a,a55808a,a55811a,a55814a,a55815a,a55818a,a55821a,a55822a,a55823a,a55826a,a55829a,a55830a,a55833a,a55837a,a55838a,a55839a,a55840a,a55843a,a55846a,a55847a,a55850a,a55853a,a55854a,a55855a,a55858a,a55861a,a55862a,a55865a,a55869a,a55870a,a55871a,a55872a,a55875a,a55878a,a55879a,a55882a,a55885a,a55886a,a55887a,a55890a,a55893a,a55894a,a55897a,a55901a,a55902a,a55903a,a55904a,a55907a,a55910a,a55911a,a55914a,a55918a,a55919a,a55920a,a55921a,a55924a,a55927a,a55928a,a55931a,a55935a,a55936a,a55937a,a55938a,a55941a,a55944a,a55945a,a55948a,a55952a,a55953a,a55954a,a55955a,a55958a,a55961a,a55962a,a55965a,a55969a,a55970a,a55971a,a55972a,a55975a,a55978a,a55979a,a55982a,a55986a,a55987a,a55988a,a55989a,a55992a,a55995a,a55996a,a55999a,a56003a,a56004a,a56005a,a56006a,a56009a,a56012a,a56013a,a56016a,a56020a,a56021a,a56022a,a56023a,a56026a,a56029a,a56030a,a56033a,a56037a,a56038a,a56039a,a56040a,a56043a,a56046a,a56047a,a56050a,a56054a,a56055a,a56056a,a56057a,a56060a,a56063a,a56064a,a56067a,a56071a,a56072a,a56073a,a56074a,a56077a,a56080a,a56081a,a56084a,a56088a,a56089a,a56090a,a56091a,a56094a,a56097a,a56098a,a56101a,a56105a,a56106a,a56107a,a56108a,a56111a,a56114a,a56115a,a56118a,a56122a,a56123a,a56124a,a56125a,a56128a,a56131a,a56132a,a56135a,a56139a,a56140a,a56141a,a56142a,a56145a,a56148a,a56149a,a56152a,a56156a,a56157a,a56158a,a56159a,a56162a,a56165a,a56166a,a56169a,a56173a,a56174a,a56175a,a56176a,a56179a,a56182a,a56183a,a56186a,a56190a,a56191a,a56192a,a56193a,a56196a,a56199a,a56200a,a56203a,a56207a,a56208a,a56209a,a56210a,a56213a,a56216a,a56217a,a56220a,a56224a,a56225a,a56226a,a56227a,a56230a,a56233a,a56234a,a56237a,a56241a,a56242a,a56243a,a56244a,a56247a,a56250a,a56251a,a56254a,a56258a,a56259a,a56260a,a56261a,a56264a,a56267a,a56268a,a56271a,a56275a,a56276a,a56277a,a56278a,a56281a,a56284a,a56285a,a56288a,a56292a,a56293a,a56294a,a56295a,a56298a,a56301a,a56302a,a56305a,a56309a,a56310a,a56311a,a56312a,a56315a,a56318a,a56319a,a56322a,a56326a,a56327a,a56328a,a56329a,a56332a,a56335a,a56336a,a56339a,a56343a,a56344a,a56345a,a56346a,a56349a,a56352a,a56353a,a56356a,a56360a,a56361a,a56362a,a56363a,a56366a,a56369a,a56370a,a56373a,a56377a,a56378a,a56379a,a56380a,a56383a,a56386a,a56387a,a56390a,a56394a,a56395a,a56396a,a56397a,a56400a,a56403a,a56404a,a56407a,a56411a,a56412a,a56413a,a56414a,a56417a,a56420a,a56421a,a56424a,a56428a,a56429a,a56430a,a56431a,a56434a,a56437a,a56438a,a56441a,a56445a,a56446a,a56447a,a56448a,a56451a,a56454a,a56455a,a56458a,a56462a,a56463a,a56464a,a56465a,a56468a,a56471a,a56472a,a56475a,a56479a,a56480a,a56481a,a56482a,a56485a,a56488a,a56489a,a56492a,a56496a,a56497a,a56498a,a56499a,a56502a,a56505a,a56506a,a56509a,a56513a,a56514a,a56515a,a56516a,a56519a,a56522a,a56523a,a56526a,a56530a,a56531a,a56532a,a56533a,a56536a,a56539a,a56540a,a56543a,a56547a,a56548a,a56549a,a56550a,a56553a,a56556a,a56557a,a56560a,a56564a,a56565a,a56566a,a56567a,a56570a,a56573a,a56574a,a56577a,a56581a,a56582a,a56583a,a56584a,a56587a,a56590a,a56591a,a56594a,a56598a,a56599a,a56600a,a56601a,a56604a,a56607a,a56608a,a56611a,a56615a,a56616a,a56617a,a56618a,a56621a,a56624a,a56625a,a56628a,a56632a,a56633a,a56634a,a56635a,a56638a,a56641a,a56642a,a56645a,a56649a,a56650a,a56651a,a56652a,a56655a,a56658a,a56659a,a56662a,a56666a,a56667a,a56668a,a56669a,a56672a,a56675a,a56676a,a56679a,a56683a,a56684a,a56685a,a56686a,a56689a,a56692a,a56693a,a56696a,a56700a,a56701a,a56702a,a56703a,a56706a,a56709a,a56710a,a56713a,a56717a,a56718a,a56719a,a56720a,a56723a,a56726a,a56727a,a56730a,a56734a,a56735a,a56736a,a56737a,a56740a,a56743a,a56744a,a56747a,a56751a,a56752a,a56753a,a56754a,a56757a,a56760a,a56761a,a56764a,a56768a,a56769a,a56770a,a56771a,a56774a,a56777a,a56778a,a56781a,a56785a,a56786a,a56787a,a56788a,a56791a,a56794a,a56795a,a56798a,a56802a,a56803a,a56804a,a56805a,a56808a,a56811a,a56812a,a56815a,a56819a,a56820a,a56821a,a56822a,a56825a,a56828a,a56829a,a56832a,a56836a,a56837a,a56838a,a56839a,a56842a,a56845a,a56846a,a56849a,a56853a,a56854a,a56855a,a56856a,a56859a,a56862a,a56863a,a56866a,a56870a,a56871a,a56872a,a56873a,a56876a,a56879a,a56880a,a56883a,a56887a,a56888a,a56889a,a56890a,a56893a,a56896a,a56897a,a56900a,a56904a,a56905a,a56906a,a56907a,a56910a,a56913a,a56914a,a56917a,a56921a,a56922a,a56923a,a56924a,a56927a,a56930a,a56931a,a56934a,a56938a,a56939a,a56940a,a56941a,a56944a,a56947a,a56948a,a56951a,a56955a,a56956a,a56957a,a56958a,a56961a,a56964a,a56965a,a56968a,a56972a,a56973a,a56974a,a56975a,a56978a,a56981a,a56982a,a56985a,a56989a,a56990a,a56991a,a56992a,a56995a,a56998a,a56999a,a57002a,a57006a,a57007a,a57008a,a57009a,a57012a,a57015a,a57016a,a57019a,a57023a,a57024a,a57025a,a57026a,a57029a,a57032a,a57033a,a57036a,a57040a,a57041a,a57042a,a57043a,a57046a,a57049a,a57050a,a57053a,a57057a,a57058a,a57059a,a57060a,a57063a,a57066a,a57067a,a57070a,a57074a,a57075a,a57076a,a57077a,a57080a,a57083a,a57084a,a57087a,a57091a,a57092a,a57093a,a57094a,a57097a,a57100a,a57101a,a57104a,a57108a,a57109a,a57110a,a57111a,a57114a,a57117a,a57118a,a57121a,a57125a,a57126a,a57127a,a57128a,a57131a,a57134a,a57135a,a57138a,a57142a,a57143a,a57144a,a57145a,a57148a,a57152a,a57153a,a57154a,a57157a,a57161a,a57162a,a57163a,a57164a,a57167a,a57170a,a57171a,a57174a,a57178a,a57179a,a57180a,a57181a,a57184a,a57188a,a57189a,a57190a,a57193a,a57197a,a57198a,a57199a,a57200a,a57203a,a57206a,a57207a,a57210a,a57214a,a57215a,a57216a,a57217a,a57220a,a57224a,a57225a,a57226a,a57229a,a57233a,a57234a,a57235a,a57236a,a57239a,a57242a,a57243a,a57246a,a57250a,a57251a,a57252a,a57253a,a57256a,a57260a,a57261a,a57262a,a57265a,a57269a,a57270a,a57271a,a57272a: std_logic;
begin

A76 <=( a6928a ) or ( a4619a );
 a1a <=( a57272a  and  a57253a );
 a2a <=( a57236a  and  a57217a );
 a3a <=( a57200a  and  a57181a );
 a4a <=( a57164a  and  a57145a );
 a5a <=( a57128a  and  a57111a );
 a6a <=( a57094a  and  a57077a );
 a7a <=( a57060a  and  a57043a );
 a8a <=( a57026a  and  a57009a );
 a9a <=( a56992a  and  a56975a );
 a10a <=( a56958a  and  a56941a );
 a11a <=( a56924a  and  a56907a );
 a12a <=( a56890a  and  a56873a );
 a13a <=( a56856a  and  a56839a );
 a14a <=( a56822a  and  a56805a );
 a15a <=( a56788a  and  a56771a );
 a16a <=( a56754a  and  a56737a );
 a17a <=( a56720a  and  a56703a );
 a18a <=( a56686a  and  a56669a );
 a19a <=( a56652a  and  a56635a );
 a20a <=( a56618a  and  a56601a );
 a21a <=( a56584a  and  a56567a );
 a22a <=( a56550a  and  a56533a );
 a23a <=( a56516a  and  a56499a );
 a24a <=( a56482a  and  a56465a );
 a25a <=( a56448a  and  a56431a );
 a26a <=( a56414a  and  a56397a );
 a27a <=( a56380a  and  a56363a );
 a28a <=( a56346a  and  a56329a );
 a29a <=( a56312a  and  a56295a );
 a30a <=( a56278a  and  a56261a );
 a31a <=( a56244a  and  a56227a );
 a32a <=( a56210a  and  a56193a );
 a33a <=( a56176a  and  a56159a );
 a34a <=( a56142a  and  a56125a );
 a35a <=( a56108a  and  a56091a );
 a36a <=( a56074a  and  a56057a );
 a37a <=( a56040a  and  a56023a );
 a38a <=( a56006a  and  a55989a );
 a39a <=( a55972a  and  a55955a );
 a40a <=( a55938a  and  a55921a );
 a41a <=( a55904a  and  a55887a );
 a42a <=( a55872a  and  a55855a );
 a43a <=( a55840a  and  a55823a );
 a44a <=( a55808a  and  a55791a );
 a45a <=( a55776a  and  a55759a );
 a46a <=( a55744a  and  a55727a );
 a47a <=( a55712a  and  a55695a );
 a48a <=( a55680a  and  a55663a );
 a49a <=( a55648a  and  a55631a );
 a50a <=( a55616a  and  a55599a );
 a51a <=( a55584a  and  a55567a );
 a52a <=( a55552a  and  a55535a );
 a53a <=( a55520a  and  a55503a );
 a54a <=( a55488a  and  a55471a );
 a55a <=( a55456a  and  a55439a );
 a56a <=( a55424a  and  a55407a );
 a57a <=( a55392a  and  a55375a );
 a58a <=( a55360a  and  a55343a );
 a59a <=( a55328a  and  a55311a );
 a60a <=( a55296a  and  a55279a );
 a61a <=( a55264a  and  a55247a );
 a62a <=( a55232a  and  a55215a );
 a63a <=( a55200a  and  a55183a );
 a64a <=( a55168a  and  a55151a );
 a65a <=( a55136a  and  a55119a );
 a66a <=( a55104a  and  a55087a );
 a67a <=( a55072a  and  a55055a );
 a68a <=( a55040a  and  a55023a );
 a69a <=( a55008a  and  a54991a );
 a70a <=( a54976a  and  a54959a );
 a71a <=( a54944a  and  a54927a );
 a72a <=( a54912a  and  a54895a );
 a73a <=( a54880a  and  a54863a );
 a74a <=( a54848a  and  a54831a );
 a75a <=( a54816a  and  a54799a );
 a76a <=( a54784a  and  a54767a );
 a77a <=( a54752a  and  a54735a );
 a78a <=( a54720a  and  a54703a );
 a79a <=( a54688a  and  a54671a );
 a80a <=( a54656a  and  a54639a );
 a81a <=( a54624a  and  a54607a );
 a82a <=( a54592a  and  a54575a );
 a83a <=( a54560a  and  a54543a );
 a84a <=( a54528a  and  a54511a );
 a85a <=( a54496a  and  a54479a );
 a86a <=( a54464a  and  a54447a );
 a87a <=( a54432a  and  a54415a );
 a88a <=( a54400a  and  a54383a );
 a89a <=( a54368a  and  a54351a );
 a90a <=( a54336a  and  a54319a );
 a91a <=( a54304a  and  a54287a );
 a92a <=( a54272a  and  a54255a );
 a93a <=( a54240a  and  a54223a );
 a94a <=( a54208a  and  a54191a );
 a95a <=( a54176a  and  a54159a );
 a96a <=( a54144a  and  a54127a );
 a97a <=( a54112a  and  a54095a );
 a98a <=( a54080a  and  a54063a );
 a99a <=( a54048a  and  a54031a );
 a100a <=( a54016a  and  a53999a );
 a101a <=( a53984a  and  a53967a );
 a102a <=( a53952a  and  a53935a );
 a103a <=( a53920a  and  a53903a );
 a104a <=( a53888a  and  a53871a );
 a105a <=( a53856a  and  a53839a );
 a106a <=( a53824a  and  a53807a );
 a107a <=( a53792a  and  a53775a );
 a108a <=( a53760a  and  a53743a );
 a109a <=( a53728a  and  a53711a );
 a110a <=( a53696a  and  a53679a );
 a111a <=( a53664a  and  a53647a );
 a112a <=( a53632a  and  a53615a );
 a113a <=( a53600a  and  a53583a );
 a114a <=( a53568a  and  a53551a );
 a115a <=( a53536a  and  a53519a );
 a116a <=( a53504a  and  a53487a );
 a117a <=( a53472a  and  a53455a );
 a118a <=( a53440a  and  a53423a );
 a119a <=( a53408a  and  a53391a );
 a120a <=( a53376a  and  a53359a );
 a121a <=( a53344a  and  a53327a );
 a122a <=( a53312a  and  a53295a );
 a123a <=( a53280a  and  a53263a );
 a124a <=( a53248a  and  a53231a );
 a125a <=( a53216a  and  a53199a );
 a126a <=( a53184a  and  a53167a );
 a127a <=( a53152a  and  a53135a );
 a128a <=( a53120a  and  a53103a );
 a129a <=( a53088a  and  a53071a );
 a130a <=( a53056a  and  a53039a );
 a131a <=( a53024a  and  a53007a );
 a132a <=( a52992a  and  a52975a );
 a133a <=( a52960a  and  a52943a );
 a134a <=( a52928a  and  a52911a );
 a135a <=( a52896a  and  a52879a );
 a136a <=( a52864a  and  a52847a );
 a137a <=( a52832a  and  a52815a );
 a138a <=( a52800a  and  a52783a );
 a139a <=( a52768a  and  a52751a );
 a140a <=( a52736a  and  a52719a );
 a141a <=( a52704a  and  a52687a );
 a142a <=( a52672a  and  a52655a );
 a143a <=( a52640a  and  a52623a );
 a144a <=( a52608a  and  a52591a );
 a145a <=( a52576a  and  a52559a );
 a146a <=( a52544a  and  a52527a );
 a147a <=( a52512a  and  a52495a );
 a148a <=( a52480a  and  a52463a );
 a149a <=( a52448a  and  a52431a );
 a150a <=( a52416a  and  a52399a );
 a151a <=( a52384a  and  a52367a );
 a152a <=( a52352a  and  a52335a );
 a153a <=( a52320a  and  a52303a );
 a154a <=( a52288a  and  a52271a );
 a155a <=( a52256a  and  a52239a );
 a156a <=( a52224a  and  a52207a );
 a157a <=( a52192a  and  a52175a );
 a158a <=( a52160a  and  a52143a );
 a159a <=( a52128a  and  a52111a );
 a160a <=( a52096a  and  a52079a );
 a161a <=( a52064a  and  a52047a );
 a162a <=( a52032a  and  a52015a );
 a163a <=( a52000a  and  a51983a );
 a164a <=( a51968a  and  a51951a );
 a165a <=( a51936a  and  a51919a );
 a166a <=( a51904a  and  a51887a );
 a167a <=( a51872a  and  a51855a );
 a168a <=( a51840a  and  a51823a );
 a169a <=( a51808a  and  a51791a );
 a170a <=( a51776a  and  a51759a );
 a171a <=( a51744a  and  a51729a );
 a172a <=( a51714a  and  a51699a );
 a173a <=( a51684a  and  a51669a );
 a174a <=( a51654a  and  a51639a );
 a175a <=( a51624a  and  a51609a );
 a176a <=( a51594a  and  a51579a );
 a177a <=( a51564a  and  a51549a );
 a178a <=( a51534a  and  a51519a );
 a179a <=( a51504a  and  a51489a );
 a180a <=( a51474a  and  a51459a );
 a181a <=( a51444a  and  a51429a );
 a182a <=( a51414a  and  a51399a );
 a183a <=( a51384a  and  a51369a );
 a184a <=( a51354a  and  a51339a );
 a185a <=( a51324a  and  a51309a );
 a186a <=( a51294a  and  a51279a );
 a187a <=( a51264a  and  a51249a );
 a188a <=( a51234a  and  a51219a );
 a189a <=( a51204a  and  a51189a );
 a190a <=( a51174a  and  a51159a );
 a191a <=( a51144a  and  a51129a );
 a192a <=( a51114a  and  a51099a );
 a193a <=( a51084a  and  a51069a );
 a194a <=( a51054a  and  a51039a );
 a195a <=( a51024a  and  a51009a );
 a196a <=( a50994a  and  a50979a );
 a197a <=( a50964a  and  a50949a );
 a198a <=( a50934a  and  a50919a );
 a199a <=( a50904a  and  a50889a );
 a200a <=( a50874a  and  a50859a );
 a201a <=( a50844a  and  a50829a );
 a202a <=( a50814a  and  a50799a );
 a203a <=( a50784a  and  a50769a );
 a204a <=( a50754a  and  a50739a );
 a205a <=( a50724a  and  a50709a );
 a206a <=( a50694a  and  a50679a );
 a207a <=( a50664a  and  a50649a );
 a208a <=( a50634a  and  a50619a );
 a209a <=( a50604a  and  a50589a );
 a210a <=( a50574a  and  a50559a );
 a211a <=( a50544a  and  a50529a );
 a212a <=( a50514a  and  a50499a );
 a213a <=( a50484a  and  a50469a );
 a214a <=( a50454a  and  a50439a );
 a215a <=( a50424a  and  a50409a );
 a216a <=( a50394a  and  a50379a );
 a217a <=( a50364a  and  a50349a );
 a218a <=( a50334a  and  a50319a );
 a219a <=( a50304a  and  a50289a );
 a220a <=( a50274a  and  a50259a );
 a221a <=( a50244a  and  a50229a );
 a222a <=( a50214a  and  a50199a );
 a223a <=( a50184a  and  a50169a );
 a224a <=( a50154a  and  a50139a );
 a225a <=( a50124a  and  a50109a );
 a226a <=( a50094a  and  a50079a );
 a227a <=( a50064a  and  a50049a );
 a228a <=( a50034a  and  a50019a );
 a229a <=( a50004a  and  a49989a );
 a230a <=( a49974a  and  a49959a );
 a231a <=( a49944a  and  a49929a );
 a232a <=( a49914a  and  a49899a );
 a233a <=( a49884a  and  a49869a );
 a234a <=( a49854a  and  a49839a );
 a235a <=( a49824a  and  a49809a );
 a236a <=( a49794a  and  a49779a );
 a237a <=( a49764a  and  a49749a );
 a238a <=( a49734a  and  a49719a );
 a239a <=( a49704a  and  a49689a );
 a240a <=( a49674a  and  a49659a );
 a241a <=( a49644a  and  a49629a );
 a242a <=( a49614a  and  a49599a );
 a243a <=( a49584a  and  a49569a );
 a244a <=( a49554a  and  a49539a );
 a245a <=( a49524a  and  a49509a );
 a246a <=( a49494a  and  a49479a );
 a247a <=( a49464a  and  a49449a );
 a248a <=( a49434a  and  a49419a );
 a249a <=( a49404a  and  a49389a );
 a250a <=( a49374a  and  a49359a );
 a251a <=( a49344a  and  a49329a );
 a252a <=( a49314a  and  a49299a );
 a253a <=( a49284a  and  a49269a );
 a254a <=( a49254a  and  a49239a );
 a255a <=( a49224a  and  a49209a );
 a256a <=( a49194a  and  a49179a );
 a257a <=( a49164a  and  a49149a );
 a258a <=( a49134a  and  a49119a );
 a259a <=( a49104a  and  a49089a );
 a260a <=( a49074a  and  a49059a );
 a261a <=( a49044a  and  a49029a );
 a262a <=( a49014a  and  a48999a );
 a263a <=( a48984a  and  a48969a );
 a264a <=( a48954a  and  a48939a );
 a265a <=( a48924a  and  a48909a );
 a266a <=( a48894a  and  a48879a );
 a267a <=( a48864a  and  a48849a );
 a268a <=( a48834a  and  a48819a );
 a269a <=( a48804a  and  a48789a );
 a270a <=( a48774a  and  a48759a );
 a271a <=( a48744a  and  a48729a );
 a272a <=( a48714a  and  a48699a );
 a273a <=( a48684a  and  a48669a );
 a274a <=( a48654a  and  a48639a );
 a275a <=( a48624a  and  a48609a );
 a276a <=( a48594a  and  a48579a );
 a277a <=( a48564a  and  a48549a );
 a278a <=( a48534a  and  a48519a );
 a279a <=( a48504a  and  a48489a );
 a280a <=( a48474a  and  a48459a );
 a281a <=( a48444a  and  a48429a );
 a282a <=( a48414a  and  a48399a );
 a283a <=( a48384a  and  a48369a );
 a284a <=( a48354a  and  a48339a );
 a285a <=( a48324a  and  a48309a );
 a286a <=( a48294a  and  a48279a );
 a287a <=( a48264a  and  a48249a );
 a288a <=( a48234a  and  a48219a );
 a289a <=( a48204a  and  a48189a );
 a290a <=( a48174a  and  a48159a );
 a291a <=( a48144a  and  a48129a );
 a292a <=( a48114a  and  a48099a );
 a293a <=( a48084a  and  a48069a );
 a294a <=( a48054a  and  a48039a );
 a295a <=( a48024a  and  a48009a );
 a296a <=( a47994a  and  a47979a );
 a297a <=( a47964a  and  a47949a );
 a298a <=( a47934a  and  a47919a );
 a299a <=( a47904a  and  a47889a );
 a300a <=( a47874a  and  a47859a );
 a301a <=( a47844a  and  a47829a );
 a302a <=( a47814a  and  a47799a );
 a303a <=( a47784a  and  a47769a );
 a304a <=( a47754a  and  a47739a );
 a305a <=( a47724a  and  a47709a );
 a306a <=( a47694a  and  a47679a );
 a307a <=( a47664a  and  a47649a );
 a308a <=( a47634a  and  a47619a );
 a309a <=( a47604a  and  a47589a );
 a310a <=( a47574a  and  a47559a );
 a311a <=( a47544a  and  a47529a );
 a312a <=( a47514a  and  a47499a );
 a313a <=( a47484a  and  a47469a );
 a314a <=( a47454a  and  a47439a );
 a315a <=( a47424a  and  a47409a );
 a316a <=( a47394a  and  a47379a );
 a317a <=( a47364a  and  a47349a );
 a318a <=( a47334a  and  a47319a );
 a319a <=( a47304a  and  a47289a );
 a320a <=( a47274a  and  a47259a );
 a321a <=( a47244a  and  a47229a );
 a322a <=( a47214a  and  a47199a );
 a323a <=( a47184a  and  a47169a );
 a324a <=( a47154a  and  a47139a );
 a325a <=( a47124a  and  a47109a );
 a326a <=( a47094a  and  a47079a );
 a327a <=( a47064a  and  a47049a );
 a328a <=( a47034a  and  a47019a );
 a329a <=( a47004a  and  a46989a );
 a330a <=( a46974a  and  a46959a );
 a331a <=( a46944a  and  a46929a );
 a332a <=( a46914a  and  a46899a );
 a333a <=( a46884a  and  a46869a );
 a334a <=( a46854a  and  a46839a );
 a335a <=( a46824a  and  a46809a );
 a336a <=( a46794a  and  a46779a );
 a337a <=( a46764a  and  a46749a );
 a338a <=( a46734a  and  a46719a );
 a339a <=( a46704a  and  a46689a );
 a340a <=( a46674a  and  a46659a );
 a341a <=( a46644a  and  a46629a );
 a342a <=( a46614a  and  a46599a );
 a343a <=( a46584a  and  a46569a );
 a344a <=( a46554a  and  a46539a );
 a345a <=( a46524a  and  a46509a );
 a346a <=( a46494a  and  a46479a );
 a347a <=( a46464a  and  a46449a );
 a348a <=( a46434a  and  a46419a );
 a349a <=( a46404a  and  a46389a );
 a350a <=( a46374a  and  a46359a );
 a351a <=( a46344a  and  a46329a );
 a352a <=( a46314a  and  a46299a );
 a353a <=( a46284a  and  a46269a );
 a354a <=( a46254a  and  a46239a );
 a355a <=( a46224a  and  a46209a );
 a356a <=( a46194a  and  a46179a );
 a357a <=( a46164a  and  a46149a );
 a358a <=( a46134a  and  a46119a );
 a359a <=( a46104a  and  a46089a );
 a360a <=( a46074a  and  a46059a );
 a361a <=( a46044a  and  a46029a );
 a362a <=( a46014a  and  a45999a );
 a363a <=( a45984a  and  a45969a );
 a364a <=( a45954a  and  a45939a );
 a365a <=( a45924a  and  a45909a );
 a366a <=( a45894a  and  a45879a );
 a367a <=( a45864a  and  a45849a );
 a368a <=( a45834a  and  a45819a );
 a369a <=( a45804a  and  a45789a );
 a370a <=( a45774a  and  a45759a );
 a371a <=( a45744a  and  a45729a );
 a372a <=( a45714a  and  a45699a );
 a373a <=( a45684a  and  a45669a );
 a374a <=( a45654a  and  a45639a );
 a375a <=( a45624a  and  a45609a );
 a376a <=( a45594a  and  a45579a );
 a377a <=( a45564a  and  a45549a );
 a378a <=( a45534a  and  a45519a );
 a379a <=( a45504a  and  a45489a );
 a380a <=( a45474a  and  a45459a );
 a381a <=( a45444a  and  a45429a );
 a382a <=( a45414a  and  a45399a );
 a383a <=( a45384a  and  a45369a );
 a384a <=( a45354a  and  a45339a );
 a385a <=( a45324a  and  a45309a );
 a386a <=( a45294a  and  a45279a );
 a387a <=( a45264a  and  a45249a );
 a388a <=( a45234a  and  a45219a );
 a389a <=( a45204a  and  a45189a );
 a390a <=( a45174a  and  a45159a );
 a391a <=( a45144a  and  a45129a );
 a392a <=( a45114a  and  a45099a );
 a393a <=( a45084a  and  a45069a );
 a394a <=( a45054a  and  a45039a );
 a395a <=( a45024a  and  a45009a );
 a396a <=( a44994a  and  a44979a );
 a397a <=( a44964a  and  a44949a );
 a398a <=( a44934a  and  a44919a );
 a399a <=( a44904a  and  a44889a );
 a400a <=( a44874a  and  a44859a );
 a401a <=( a44844a  and  a44829a );
 a402a <=( a44814a  and  a44799a );
 a403a <=( a44784a  and  a44769a );
 a404a <=( a44754a  and  a44739a );
 a405a <=( a44724a  and  a44709a );
 a406a <=( a44694a  and  a44679a );
 a407a <=( a44664a  and  a44649a );
 a408a <=( a44634a  and  a44619a );
 a409a <=( a44604a  and  a44589a );
 a410a <=( a44574a  and  a44559a );
 a411a <=( a44544a  and  a44529a );
 a412a <=( a44516a  and  a44501a );
 a413a <=( a44488a  and  a44473a );
 a414a <=( a44460a  and  a44445a );
 a415a <=( a44432a  and  a44417a );
 a416a <=( a44404a  and  a44389a );
 a417a <=( a44376a  and  a44361a );
 a418a <=( a44348a  and  a44333a );
 a419a <=( a44320a  and  a44305a );
 a420a <=( a44292a  and  a44277a );
 a421a <=( a44264a  and  a44249a );
 a422a <=( a44236a  and  a44221a );
 a423a <=( a44208a  and  a44193a );
 a424a <=( a44180a  and  a44165a );
 a425a <=( a44152a  and  a44137a );
 a426a <=( a44124a  and  a44109a );
 a427a <=( a44096a  and  a44081a );
 a428a <=( a44068a  and  a44053a );
 a429a <=( a44040a  and  a44025a );
 a430a <=( a44012a  and  a43997a );
 a431a <=( a43984a  and  a43969a );
 a432a <=( a43956a  and  a43941a );
 a433a <=( a43928a  and  a43913a );
 a434a <=( a43900a  and  a43885a );
 a435a <=( a43872a  and  a43857a );
 a436a <=( a43844a  and  a43829a );
 a437a <=( a43816a  and  a43801a );
 a438a <=( a43788a  and  a43773a );
 a439a <=( a43760a  and  a43745a );
 a440a <=( a43732a  and  a43717a );
 a441a <=( a43704a  and  a43689a );
 a442a <=( a43676a  and  a43661a );
 a443a <=( a43648a  and  a43633a );
 a444a <=( a43620a  and  a43605a );
 a445a <=( a43592a  and  a43577a );
 a446a <=( a43564a  and  a43549a );
 a447a <=( a43536a  and  a43521a );
 a448a <=( a43508a  and  a43493a );
 a449a <=( a43480a  and  a43465a );
 a450a <=( a43452a  and  a43437a );
 a451a <=( a43424a  and  a43409a );
 a452a <=( a43396a  and  a43381a );
 a453a <=( a43368a  and  a43353a );
 a454a <=( a43340a  and  a43325a );
 a455a <=( a43312a  and  a43297a );
 a456a <=( a43284a  and  a43269a );
 a457a <=( a43256a  and  a43241a );
 a458a <=( a43228a  and  a43213a );
 a459a <=( a43200a  and  a43185a );
 a460a <=( a43172a  and  a43157a );
 a461a <=( a43144a  and  a43129a );
 a462a <=( a43116a  and  a43101a );
 a463a <=( a43088a  and  a43073a );
 a464a <=( a43060a  and  a43045a );
 a465a <=( a43032a  and  a43017a );
 a466a <=( a43004a  and  a42989a );
 a467a <=( a42976a  and  a42961a );
 a468a <=( a42948a  and  a42933a );
 a469a <=( a42920a  and  a42905a );
 a470a <=( a42892a  and  a42877a );
 a471a <=( a42864a  and  a42849a );
 a472a <=( a42836a  and  a42821a );
 a473a <=( a42808a  and  a42793a );
 a474a <=( a42780a  and  a42765a );
 a475a <=( a42752a  and  a42737a );
 a476a <=( a42724a  and  a42709a );
 a477a <=( a42696a  and  a42681a );
 a478a <=( a42668a  and  a42653a );
 a479a <=( a42640a  and  a42625a );
 a480a <=( a42612a  and  a42597a );
 a481a <=( a42584a  and  a42569a );
 a482a <=( a42556a  and  a42541a );
 a483a <=( a42528a  and  a42513a );
 a484a <=( a42500a  and  a42485a );
 a485a <=( a42472a  and  a42457a );
 a486a <=( a42444a  and  a42429a );
 a487a <=( a42416a  and  a42401a );
 a488a <=( a42388a  and  a42373a );
 a489a <=( a42360a  and  a42345a );
 a490a <=( a42332a  and  a42317a );
 a491a <=( a42304a  and  a42289a );
 a492a <=( a42276a  and  a42261a );
 a493a <=( a42248a  and  a42233a );
 a494a <=( a42220a  and  a42205a );
 a495a <=( a42192a  and  a42177a );
 a496a <=( a42164a  and  a42149a );
 a497a <=( a42136a  and  a42121a );
 a498a <=( a42108a  and  a42093a );
 a499a <=( a42080a  and  a42065a );
 a500a <=( a42052a  and  a42037a );
 a501a <=( a42024a  and  a42009a );
 a502a <=( a41996a  and  a41981a );
 a503a <=( a41968a  and  a41953a );
 a504a <=( a41940a  and  a41925a );
 a505a <=( a41912a  and  a41897a );
 a506a <=( a41884a  and  a41869a );
 a507a <=( a41856a  and  a41841a );
 a508a <=( a41828a  and  a41813a );
 a509a <=( a41800a  and  a41785a );
 a510a <=( a41772a  and  a41757a );
 a511a <=( a41744a  and  a41729a );
 a512a <=( a41716a  and  a41701a );
 a513a <=( a41688a  and  a41673a );
 a514a <=( a41660a  and  a41645a );
 a515a <=( a41632a  and  a41617a );
 a516a <=( a41604a  and  a41589a );
 a517a <=( a41576a  and  a41561a );
 a518a <=( a41548a  and  a41533a );
 a519a <=( a41520a  and  a41505a );
 a520a <=( a41492a  and  a41477a );
 a521a <=( a41464a  and  a41449a );
 a522a <=( a41436a  and  a41421a );
 a523a <=( a41408a  and  a41393a );
 a524a <=( a41380a  and  a41365a );
 a525a <=( a41352a  and  a41337a );
 a526a <=( a41324a  and  a41309a );
 a527a <=( a41296a  and  a41281a );
 a528a <=( a41268a  and  a41253a );
 a529a <=( a41240a  and  a41225a );
 a530a <=( a41212a  and  a41197a );
 a531a <=( a41184a  and  a41169a );
 a532a <=( a41156a  and  a41141a );
 a533a <=( a41128a  and  a41113a );
 a534a <=( a41100a  and  a41085a );
 a535a <=( a41072a  and  a41057a );
 a536a <=( a41044a  and  a41029a );
 a537a <=( a41016a  and  a41001a );
 a538a <=( a40988a  and  a40973a );
 a539a <=( a40960a  and  a40945a );
 a540a <=( a40932a  and  a40917a );
 a541a <=( a40904a  and  a40889a );
 a542a <=( a40876a  and  a40861a );
 a543a <=( a40848a  and  a40833a );
 a544a <=( a40820a  and  a40805a );
 a545a <=( a40792a  and  a40777a );
 a546a <=( a40764a  and  a40749a );
 a547a <=( a40736a  and  a40721a );
 a548a <=( a40708a  and  a40693a );
 a549a <=( a40680a  and  a40665a );
 a550a <=( a40652a  and  a40637a );
 a551a <=( a40624a  and  a40609a );
 a552a <=( a40596a  and  a40581a );
 a553a <=( a40568a  and  a40553a );
 a554a <=( a40540a  and  a40525a );
 a555a <=( a40512a  and  a40497a );
 a556a <=( a40484a  and  a40469a );
 a557a <=( a40456a  and  a40441a );
 a558a <=( a40428a  and  a40413a );
 a559a <=( a40400a  and  a40385a );
 a560a <=( a40372a  and  a40357a );
 a561a <=( a40344a  and  a40329a );
 a562a <=( a40316a  and  a40301a );
 a563a <=( a40288a  and  a40273a );
 a564a <=( a40260a  and  a40245a );
 a565a <=( a40232a  and  a40217a );
 a566a <=( a40204a  and  a40189a );
 a567a <=( a40176a  and  a40161a );
 a568a <=( a40148a  and  a40133a );
 a569a <=( a40120a  and  a40105a );
 a570a <=( a40092a  and  a40077a );
 a571a <=( a40064a  and  a40049a );
 a572a <=( a40036a  and  a40021a );
 a573a <=( a40008a  and  a39993a );
 a574a <=( a39980a  and  a39965a );
 a575a <=( a39952a  and  a39937a );
 a576a <=( a39924a  and  a39909a );
 a577a <=( a39896a  and  a39881a );
 a578a <=( a39868a  and  a39853a );
 a579a <=( a39840a  and  a39825a );
 a580a <=( a39812a  and  a39797a );
 a581a <=( a39784a  and  a39769a );
 a582a <=( a39756a  and  a39741a );
 a583a <=( a39728a  and  a39713a );
 a584a <=( a39700a  and  a39685a );
 a585a <=( a39672a  and  a39657a );
 a586a <=( a39644a  and  a39629a );
 a587a <=( a39616a  and  a39601a );
 a588a <=( a39588a  and  a39573a );
 a589a <=( a39560a  and  a39545a );
 a590a <=( a39532a  and  a39517a );
 a591a <=( a39504a  and  a39489a );
 a592a <=( a39476a  and  a39461a );
 a593a <=( a39448a  and  a39433a );
 a594a <=( a39420a  and  a39405a );
 a595a <=( a39392a  and  a39377a );
 a596a <=( a39364a  and  a39349a );
 a597a <=( a39336a  and  a39321a );
 a598a <=( a39308a  and  a39293a );
 a599a <=( a39280a  and  a39265a );
 a600a <=( a39252a  and  a39237a );
 a601a <=( a39224a  and  a39209a );
 a602a <=( a39196a  and  a39181a );
 a603a <=( a39168a  and  a39153a );
 a604a <=( a39140a  and  a39125a );
 a605a <=( a39112a  and  a39097a );
 a606a <=( a39084a  and  a39069a );
 a607a <=( a39056a  and  a39041a );
 a608a <=( a39028a  and  a39013a );
 a609a <=( a39000a  and  a38985a );
 a610a <=( a38972a  and  a38957a );
 a611a <=( a38944a  and  a38929a );
 a612a <=( a38916a  and  a38901a );
 a613a <=( a38888a  and  a38873a );
 a614a <=( a38860a  and  a38845a );
 a615a <=( a38832a  and  a38817a );
 a616a <=( a38804a  and  a38789a );
 a617a <=( a38776a  and  a38761a );
 a618a <=( a38748a  and  a38733a );
 a619a <=( a38720a  and  a38705a );
 a620a <=( a38692a  and  a38677a );
 a621a <=( a38664a  and  a38649a );
 a622a <=( a38636a  and  a38621a );
 a623a <=( a38608a  and  a38593a );
 a624a <=( a38580a  and  a38565a );
 a625a <=( a38552a  and  a38537a );
 a626a <=( a38524a  and  a38509a );
 a627a <=( a38496a  and  a38481a );
 a628a <=( a38468a  and  a38453a );
 a629a <=( a38440a  and  a38425a );
 a630a <=( a38412a  and  a38397a );
 a631a <=( a38384a  and  a38369a );
 a632a <=( a38356a  and  a38341a );
 a633a <=( a38328a  and  a38313a );
 a634a <=( a38300a  and  a38285a );
 a635a <=( a38272a  and  a38257a );
 a636a <=( a38244a  and  a38229a );
 a637a <=( a38216a  and  a38201a );
 a638a <=( a38188a  and  a38173a );
 a639a <=( a38160a  and  a38145a );
 a640a <=( a38132a  and  a38117a );
 a641a <=( a38104a  and  a38089a );
 a642a <=( a38076a  and  a38061a );
 a643a <=( a38048a  and  a38033a );
 a644a <=( a38020a  and  a38005a );
 a645a <=( a37992a  and  a37977a );
 a646a <=( a37964a  and  a37949a );
 a647a <=( a37936a  and  a37921a );
 a648a <=( a37908a  and  a37893a );
 a649a <=( a37880a  and  a37865a );
 a650a <=( a37852a  and  a37837a );
 a651a <=( a37824a  and  a37811a );
 a652a <=( a37798a  and  a37785a );
 a653a <=( a37772a  and  a37759a );
 a654a <=( a37746a  and  a37733a );
 a655a <=( a37720a  and  a37707a );
 a656a <=( a37694a  and  a37681a );
 a657a <=( a37668a  and  a37655a );
 a658a <=( a37642a  and  a37629a );
 a659a <=( a37616a  and  a37603a );
 a660a <=( a37590a  and  a37577a );
 a661a <=( a37564a  and  a37551a );
 a662a <=( a37538a  and  a37525a );
 a663a <=( a37512a  and  a37499a );
 a664a <=( a37486a  and  a37473a );
 a665a <=( a37460a  and  a37447a );
 a666a <=( a37434a  and  a37421a );
 a667a <=( a37408a  and  a37395a );
 a668a <=( a37382a  and  a37369a );
 a669a <=( a37356a  and  a37343a );
 a670a <=( a37330a  and  a37317a );
 a671a <=( a37304a  and  a37291a );
 a672a <=( a37278a  and  a37265a );
 a673a <=( a37252a  and  a37239a );
 a674a <=( a37226a  and  a37213a );
 a675a <=( a37200a  and  a37187a );
 a676a <=( a37174a  and  a37161a );
 a677a <=( a37148a  and  a37135a );
 a678a <=( a37122a  and  a37109a );
 a679a <=( a37096a  and  a37083a );
 a680a <=( a37070a  and  a37057a );
 a681a <=( a37044a  and  a37031a );
 a682a <=( a37018a  and  a37005a );
 a683a <=( a36992a  and  a36979a );
 a684a <=( a36966a  and  a36953a );
 a685a <=( a36940a  and  a36927a );
 a686a <=( a36914a  and  a36901a );
 a687a <=( a36888a  and  a36875a );
 a688a <=( a36862a  and  a36849a );
 a689a <=( a36836a  and  a36823a );
 a690a <=( a36810a  and  a36797a );
 a691a <=( a36784a  and  a36771a );
 a692a <=( a36758a  and  a36745a );
 a693a <=( a36732a  and  a36719a );
 a694a <=( a36706a  and  a36693a );
 a695a <=( a36680a  and  a36667a );
 a696a <=( a36654a  and  a36641a );
 a697a <=( a36628a  and  a36615a );
 a698a <=( a36602a  and  a36589a );
 a699a <=( a36576a  and  a36563a );
 a700a <=( a36550a  and  a36537a );
 a701a <=( a36524a  and  a36511a );
 a702a <=( a36498a  and  a36485a );
 a703a <=( a36472a  and  a36459a );
 a704a <=( a36446a  and  a36433a );
 a705a <=( a36420a  and  a36407a );
 a706a <=( a36394a  and  a36381a );
 a707a <=( a36368a  and  a36355a );
 a708a <=( a36342a  and  a36329a );
 a709a <=( a36316a  and  a36303a );
 a710a <=( a36290a  and  a36277a );
 a711a <=( a36264a  and  a36251a );
 a712a <=( a36238a  and  a36225a );
 a713a <=( a36212a  and  a36199a );
 a714a <=( a36186a  and  a36173a );
 a715a <=( a36160a  and  a36147a );
 a716a <=( a36134a  and  a36121a );
 a717a <=( a36108a  and  a36095a );
 a718a <=( a36082a  and  a36069a );
 a719a <=( a36056a  and  a36043a );
 a720a <=( a36030a  and  a36017a );
 a721a <=( a36004a  and  a35991a );
 a722a <=( a35978a  and  a35965a );
 a723a <=( a35952a  and  a35939a );
 a724a <=( a35926a  and  a35913a );
 a725a <=( a35900a  and  a35887a );
 a726a <=( a35874a  and  a35861a );
 a727a <=( a35848a  and  a35835a );
 a728a <=( a35822a  and  a35809a );
 a729a <=( a35796a  and  a35783a );
 a730a <=( a35770a  and  a35757a );
 a731a <=( a35744a  and  a35731a );
 a732a <=( a35718a  and  a35705a );
 a733a <=( a35692a  and  a35679a );
 a734a <=( a35666a  and  a35653a );
 a735a <=( a35640a  and  a35627a );
 a736a <=( a35614a  and  a35601a );
 a737a <=( a35588a  and  a35575a );
 a738a <=( a35562a  and  a35549a );
 a739a <=( a35536a  and  a35523a );
 a740a <=( a35510a  and  a35497a );
 a741a <=( a35484a  and  a35471a );
 a742a <=( a35458a  and  a35445a );
 a743a <=( a35432a  and  a35419a );
 a744a <=( a35406a  and  a35393a );
 a745a <=( a35380a  and  a35367a );
 a746a <=( a35354a  and  a35341a );
 a747a <=( a35328a  and  a35315a );
 a748a <=( a35302a  and  a35289a );
 a749a <=( a35276a  and  a35263a );
 a750a <=( a35250a  and  a35237a );
 a751a <=( a35224a  and  a35211a );
 a752a <=( a35198a  and  a35185a );
 a753a <=( a35172a  and  a35159a );
 a754a <=( a35146a  and  a35133a );
 a755a <=( a35120a  and  a35107a );
 a756a <=( a35094a  and  a35081a );
 a757a <=( a35068a  and  a35055a );
 a758a <=( a35042a  and  a35029a );
 a759a <=( a35016a  and  a35003a );
 a760a <=( a34990a  and  a34977a );
 a761a <=( a34964a  and  a34951a );
 a762a <=( a34938a  and  a34925a );
 a763a <=( a34912a  and  a34899a );
 a764a <=( a34886a  and  a34873a );
 a765a <=( a34860a  and  a34847a );
 a766a <=( a34834a  and  a34821a );
 a767a <=( a34808a  and  a34795a );
 a768a <=( a34782a  and  a34769a );
 a769a <=( a34756a  and  a34743a );
 a770a <=( a34730a  and  a34717a );
 a771a <=( a34704a  and  a34691a );
 a772a <=( a34678a  and  a34665a );
 a773a <=( a34652a  and  a34639a );
 a774a <=( a34626a  and  a34613a );
 a775a <=( a34600a  and  a34587a );
 a776a <=( a34574a  and  a34561a );
 a777a <=( a34548a  and  a34535a );
 a778a <=( a34522a  and  a34509a );
 a779a <=( a34496a  and  a34483a );
 a780a <=( a34472a  and  a34459a );
 a781a <=( a34448a  and  a34435a );
 a782a <=( a34424a  and  a34411a );
 a783a <=( a34400a  and  a34387a );
 a784a <=( a34376a  and  a34363a );
 a785a <=( a34352a  and  a34339a );
 a786a <=( a34328a  and  a34315a );
 a787a <=( a34304a  and  a34291a );
 a788a <=( a34280a  and  a34267a );
 a789a <=( a34256a  and  a34243a );
 a790a <=( a34232a  and  a34219a );
 a791a <=( a34208a  and  a34195a );
 a792a <=( a34184a  and  a34171a );
 a793a <=( a34160a  and  a34147a );
 a794a <=( a34136a  and  a34123a );
 a795a <=( a34112a  and  a34099a );
 a796a <=( a34088a  and  a34075a );
 a797a <=( a34064a  and  a34051a );
 a798a <=( a34040a  and  a34027a );
 a799a <=( a34016a  and  a34003a );
 a800a <=( a33992a  and  a33979a );
 a801a <=( a33968a  and  a33955a );
 a802a <=( a33944a  and  a33931a );
 a803a <=( a33920a  and  a33907a );
 a804a <=( a33896a  and  a33883a );
 a805a <=( a33872a  and  a33859a );
 a806a <=( a33848a  and  a33835a );
 a807a <=( a33824a  and  a33811a );
 a808a <=( a33800a  and  a33787a );
 a809a <=( a33776a  and  a33763a );
 a810a <=( a33752a  and  a33739a );
 a811a <=( a33728a  and  a33715a );
 a812a <=( a33704a  and  a33691a );
 a813a <=( a33680a  and  a33667a );
 a814a <=( a33656a  and  a33643a );
 a815a <=( a33632a  and  a33619a );
 a816a <=( a33608a  and  a33595a );
 a817a <=( a33584a  and  a33571a );
 a818a <=( a33560a  and  a33547a );
 a819a <=( a33536a  and  a33523a );
 a820a <=( a33512a  and  a33499a );
 a821a <=( a33488a  and  a33475a );
 a822a <=( a33464a  and  a33451a );
 a823a <=( a33440a  and  a33427a );
 a824a <=( a33416a  and  a33403a );
 a825a <=( a33392a  and  a33379a );
 a826a <=( a33368a  and  a33355a );
 a827a <=( a33344a  and  a33331a );
 a828a <=( a33320a  and  a33307a );
 a829a <=( a33296a  and  a33283a );
 a830a <=( a33272a  and  a33259a );
 a831a <=( a33248a  and  a33235a );
 a832a <=( a33224a  and  a33211a );
 a833a <=( a33200a  and  a33187a );
 a834a <=( a33176a  and  a33163a );
 a835a <=( a33152a  and  a33139a );
 a836a <=( a33128a  and  a33115a );
 a837a <=( a33104a  and  a33091a );
 a838a <=( a33080a  and  a33067a );
 a839a <=( a33056a  and  a33043a );
 a840a <=( a33032a  and  a33019a );
 a841a <=( a33008a  and  a32995a );
 a842a <=( a32984a  and  a32971a );
 a843a <=( a32960a  and  a32949a );
 a844a <=( a32938a  and  a32927a );
 a845a <=( a32916a  and  a32905a );
 a846a <=( a32894a  and  a32883a );
 a847a <=( a32872a  and  a32861a );
 a848a <=( a32850a  and  a32839a );
 a849a <=( a32828a  and  a32817a );
 a850a <=( a32806a  and  a32795a );
 a851a <=( a32784a  and  a32773a );
 a852a <=( a32762a  and  a32751a );
 a853a <=( a32740a  and  a32729a );
 a854a <=( a32718a  and  a32707a );
 a855a <=( a32696a  and  a32685a );
 a856a <=( a32674a  and  a32663a );
 a857a <=( a32652a  and  a32641a );
 a858a <=( a32630a  and  a32619a );
 a859a <=( a32608a  and  a32597a );
 a860a <=( a32586a  and  a32575a );
 a861a <=( a32564a  and  a32553a );
 a862a <=( a32542a  and  a32531a );
 a863a <=( a32520a  and  a32509a );
 a864a <=( a32498a  and  a32487a );
 a865a <=( a32476a  and  a32465a );
 a866a <=( a32454a  and  a32443a );
 a867a <=( a32432a  and  a32421a );
 a868a <=( a32410a  and  a32399a );
 a869a <=( a32388a  and  a32377a );
 a870a <=( a32366a  and  a32355a );
 a871a <=( a32344a  and  a32333a );
 a872a <=( a32322a  and  a32311a );
 a873a <=( a32300a  and  a32289a );
 a874a <=( a32278a  and  a32267a );
 a875a <=( a32256a  and  a32245a );
 a876a <=( a32234a  and  a32223a );
 a877a <=( a32212a  and  a32201a );
 a878a <=( a32190a  and  a32179a );
 a879a <=( a32168a  and  a32157a );
 a880a <=( a32146a  and  a32135a );
 a881a <=( a32124a  and  a32113a );
 a882a <=( a32102a  and  a32091a );
 a883a <=( a32080a  and  a32069a );
 a884a <=( a32058a  and  a32047a );
 a885a <=( a32036a  and  a32025a );
 a886a <=( a32014a  and  a32003a );
 a887a <=( a31992a  and  a31981a );
 a888a <=( a31970a  and  a31959a );
 a889a <=( a31948a  and  a31937a );
 a890a <=( a31926a  and  a31915a );
 a891a <=( a31904a  and  a31893a );
 a892a <=( a31882a  and  a31871a );
 a893a <=( a31860a  and  a31849a );
 a894a <=( a31838a  and  a31827a );
 a895a <=( a31816a  and  a31805a );
 a896a <=( a31794a  and  a31783a );
 a897a <=( a31772a  and  a31761a );
 a898a <=( a31750a  and  a31739a );
 a899a <=( a31728a  and  a31717a );
 a900a <=( a31706a  and  a31695a );
 a901a <=( a31684a  and  a31673a );
 a902a <=( a31662a  and  a31651a );
 a903a <=( a31640a  and  a31629a );
 a904a <=( a31618a  and  a31607a );
 a905a <=( a31596a  and  a31585a );
 a906a <=( a31574a  and  a31563a );
 a907a <=( a31552a  and  a31541a );
 a908a <=( a31530a  and  a31519a );
 a909a <=( a31508a  and  a31497a );
 a910a <=( a31486a  and  a31475a );
 a911a <=( a31464a  and  a31453a );
 a912a <=( a31442a  and  a31431a );
 a913a <=( a31420a  and  a31409a );
 a914a <=( a31398a  and  a31387a );
 a915a <=( a31376a  and  a31365a );
 a916a <=( a31354a  and  a31343a );
 a917a <=( a31332a  and  a31321a );
 a918a <=( a31310a  and  a31299a );
 a919a <=( a31288a  and  a31277a );
 a920a <=( a31266a  and  a31255a );
 a921a <=( a31244a  and  a31233a );
 a922a <=( a31222a  and  a31211a );
 a923a <=( a31200a  and  a31189a );
 a924a <=( a31178a  and  a31167a );
 a925a <=( a31156a  and  a31145a );
 a926a <=( a31134a  and  a31123a );
 a927a <=( a31112a  and  a31101a );
 a928a <=( a31090a  and  a31079a );
 a929a <=( a31068a  and  a31057a );
 a930a <=( a31046a  and  a31035a );
 a931a <=( a31024a  and  a31013a );
 a932a <=( a31002a  and  a30991a );
 a933a <=( a30980a  and  a30969a );
 a934a <=( a30958a  and  a30947a );
 a935a <=( a30936a  and  a30925a );
 a936a <=( a30914a  and  a30903a );
 a937a <=( a30892a  and  a30881a );
 a938a <=( a30870a  and  a30859a );
 a939a <=( a30848a  and  a30837a );
 a940a <=( a30826a  and  a30815a );
 a941a <=( a30804a  and  a30793a );
 a942a <=( a30782a  and  a30771a );
 a943a <=( a30760a  and  a30749a );
 a944a <=( a30738a  and  a30727a );
 a945a <=( a30716a  and  a30705a );
 a946a <=( a30694a  and  a30683a );
 a947a <=( a30672a  and  a30661a );
 a948a <=( a30650a  and  a30639a );
 a949a <=( a30628a  and  a30617a );
 a950a <=( a30606a  and  a30595a );
 a951a <=( a30584a  and  a30573a );
 a952a <=( a30562a  and  a30551a );
 a953a <=( a30540a  and  a30529a );
 a954a <=( a30518a  and  a30507a );
 a955a <=( a30496a  and  a30485a );
 a956a <=( a30474a  and  a30463a );
 a957a <=( a30452a  and  a30441a );
 a958a <=( a30430a  and  a30419a );
 a959a <=( a30408a  and  a30397a );
 a960a <=( a30386a  and  a30375a );
 a961a <=( a30364a  and  a30353a );
 a962a <=( a30342a  and  a30331a );
 a963a <=( a30320a  and  a30309a );
 a964a <=( a30298a  and  a30287a );
 a965a <=( a30276a  and  a30265a );
 a966a <=( a30254a  and  a30243a );
 a967a <=( a30232a  and  a30221a );
 a968a <=( a30210a  and  a30199a );
 a969a <=( a30188a  and  a30177a );
 a970a <=( a30166a  and  a30155a );
 a971a <=( a30144a  and  a30133a );
 a972a <=( a30122a  and  a30111a );
 a973a <=( a30100a  and  a30089a );
 a974a <=( a30078a  and  a30067a );
 a975a <=( a30056a  and  a30045a );
 a976a <=( a30034a  and  a30023a );
 a977a <=( a30012a  and  a30001a );
 a978a <=( a29990a  and  a29979a );
 a979a <=( a29968a  and  a29957a );
 a980a <=( a29946a  and  a29935a );
 a981a <=( a29924a  and  a29913a );
 a982a <=( a29902a  and  a29891a );
 a983a <=( a29880a  and  a29869a );
 a984a <=( a29858a  and  a29847a );
 a985a <=( a29836a  and  a29825a );
 a986a <=( a29814a  and  a29803a );
 a987a <=( a29792a  and  a29781a );
 a988a <=( a29770a  and  a29759a );
 a989a <=( a29748a  and  a29737a );
 a990a <=( a29726a  and  a29715a );
 a991a <=( a29704a  and  a29693a );
 a992a <=( a29682a  and  a29671a );
 a993a <=( a29660a  and  a29649a );
 a994a <=( a29638a  and  a29627a );
 a995a <=( a29616a  and  a29605a );
 a996a <=( a29594a  and  a29583a );
 a997a <=( a29572a  and  a29561a );
 a998a <=( a29550a  and  a29539a );
 a999a <=( a29528a  and  a29517a );
 a1000a <=( a29506a  and  a29495a );
 a1001a <=( a29484a  and  a29473a );
 a1002a <=( a29462a  and  a29451a );
 a1003a <=( a29440a  and  a29429a );
 a1004a <=( a29420a  and  a29409a );
 a1005a <=( a29400a  and  a29389a );
 a1006a <=( a29380a  and  a29369a );
 a1007a <=( a29360a  and  a29349a );
 a1008a <=( a29340a  and  a29329a );
 a1009a <=( a29320a  and  a29309a );
 a1010a <=( a29300a  and  a29289a );
 a1011a <=( a29280a  and  a29269a );
 a1012a <=( a29260a  and  a29249a );
 a1013a <=( a29240a  and  a29229a );
 a1014a <=( a29220a  and  a29209a );
 a1015a <=( a29200a  and  a29189a );
 a1016a <=( a29180a  and  a29169a );
 a1017a <=( a29160a  and  a29149a );
 a1018a <=( a29140a  and  a29129a );
 a1019a <=( a29120a  and  a29109a );
 a1020a <=( a29100a  and  a29089a );
 a1021a <=( a29080a  and  a29069a );
 a1022a <=( a29060a  and  a29049a );
 a1023a <=( a29040a  and  a29029a );
 a1024a <=( a29020a  and  a29009a );
 a1025a <=( a29000a  and  a28989a );
 a1026a <=( a28980a  and  a28969a );
 a1027a <=( a28960a  and  a28949a );
 a1028a <=( a28940a  and  a28929a );
 a1029a <=( a28920a  and  a28909a );
 a1030a <=( a28900a  and  a28889a );
 a1031a <=( a28880a  and  a28869a );
 a1032a <=( a28860a  and  a28849a );
 a1033a <=( a28840a  and  a28829a );
 a1034a <=( a28820a  and  a28809a );
 a1035a <=( a28800a  and  a28789a );
 a1036a <=( a28780a  and  a28769a );
 a1037a <=( a28760a  and  a28749a );
 a1038a <=( a28740a  and  a28729a );
 a1039a <=( a28720a  and  a28709a );
 a1040a <=( a28700a  and  a28689a );
 a1041a <=( a28680a  and  a28669a );
 a1042a <=( a28660a  and  a28649a );
 a1043a <=( a28640a  and  a28629a );
 a1044a <=( a28620a  and  a28609a );
 a1045a <=( a28600a  and  a28589a );
 a1046a <=( a28580a  and  a28569a );
 a1047a <=( a28560a  and  a28549a );
 a1048a <=( a28540a  and  a28529a );
 a1049a <=( a28520a  and  a28509a );
 a1050a <=( a28500a  and  a28489a );
 a1051a <=( a28480a  and  a28469a );
 a1052a <=( a28460a  and  a28449a );
 a1053a <=( a28440a  and  a28429a );
 a1054a <=( a28420a  and  a28409a );
 a1055a <=( a28400a  and  a28389a );
 a1056a <=( a28380a  and  a28369a );
 a1057a <=( a28360a  and  a28349a );
 a1058a <=( a28340a  and  a28329a );
 a1059a <=( a28320a  and  a28309a );
 a1060a <=( a28300a  and  a28289a );
 a1061a <=( a28280a  and  a28269a );
 a1062a <=( a28260a  and  a28249a );
 a1063a <=( a28240a  and  a28229a );
 a1064a <=( a28220a  and  a28209a );
 a1065a <=( a28200a  and  a28189a );
 a1066a <=( a28180a  and  a28169a );
 a1067a <=( a28160a  and  a28149a );
 a1068a <=( a28140a  and  a28129a );
 a1069a <=( a28120a  and  a28109a );
 a1070a <=( a28100a  and  a28089a );
 a1071a <=( a28080a  and  a28069a );
 a1072a <=( a28060a  and  a28049a );
 a1073a <=( a28040a  and  a28029a );
 a1074a <=( a28020a  and  a28009a );
 a1075a <=( a28000a  and  a27989a );
 a1076a <=( a27980a  and  a27969a );
 a1077a <=( a27960a  and  a27949a );
 a1078a <=( a27940a  and  a27929a );
 a1079a <=( a27920a  and  a27909a );
 a1080a <=( a27900a  and  a27889a );
 a1081a <=( a27880a  and  a27869a );
 a1082a <=( a27860a  and  a27849a );
 a1083a <=( a27840a  and  a27829a );
 a1084a <=( a27820a  and  a27809a );
 a1085a <=( a27800a  and  a27789a );
 a1086a <=( a27780a  and  a27769a );
 a1087a <=( a27760a  and  a27749a );
 a1088a <=( a27740a  and  a27729a );
 a1089a <=( a27720a  and  a27709a );
 a1090a <=( a27700a  and  a27689a );
 a1091a <=( a27680a  and  a27669a );
 a1092a <=( a27660a  and  a27649a );
 a1093a <=( a27640a  and  a27629a );
 a1094a <=( a27620a  and  a27609a );
 a1095a <=( a27600a  and  a27589a );
 a1096a <=( a27580a  and  a27569a );
 a1097a <=( a27560a  and  a27549a );
 a1098a <=( a27540a  and  a27529a );
 a1099a <=( a27520a  and  a27509a );
 a1100a <=( a27500a  and  a27489a );
 a1101a <=( a27480a  and  a27469a );
 a1102a <=( a27460a  and  a27449a );
 a1103a <=( a27440a  and  a27429a );
 a1104a <=( a27420a  and  a27409a );
 a1105a <=( a27400a  and  a27389a );
 a1106a <=( a27380a  and  a27369a );
 a1107a <=( a27360a  and  a27349a );
 a1108a <=( a27340a  and  a27329a );
 a1109a <=( a27320a  and  a27309a );
 a1110a <=( a27300a  and  a27289a );
 a1111a <=( a27280a  and  a27269a );
 a1112a <=( a27260a  and  a27249a );
 a1113a <=( a27240a  and  a27229a );
 a1114a <=( a27220a  and  a27209a );
 a1115a <=( a27200a  and  a27189a );
 a1116a <=( a27180a  and  a27169a );
 a1117a <=( a27160a  and  a27149a );
 a1118a <=( a27140a  and  a27129a );
 a1119a <=( a27120a  and  a27109a );
 a1120a <=( a27100a  and  a27089a );
 a1121a <=( a27080a  and  a27069a );
 a1122a <=( a27060a  and  a27049a );
 a1123a <=( a27040a  and  a27029a );
 a1124a <=( a27020a  and  a27009a );
 a1125a <=( a27000a  and  a26989a );
 a1126a <=( a26980a  and  a26969a );
 a1127a <=( a26960a  and  a26949a );
 a1128a <=( a26940a  and  a26929a );
 a1129a <=( a26920a  and  a26909a );
 a1130a <=( a26900a  and  a26889a );
 a1131a <=( a26880a  and  a26869a );
 a1132a <=( a26860a  and  a26849a );
 a1133a <=( a26840a  and  a26829a );
 a1134a <=( a26820a  and  a26809a );
 a1135a <=( a26800a  and  a26789a );
 a1136a <=( a26780a  and  a26769a );
 a1137a <=( a26760a  and  a26749a );
 a1138a <=( a26740a  and  a26729a );
 a1139a <=( a26720a  and  a26709a );
 a1140a <=( a26700a  and  a26689a );
 a1141a <=( a26680a  and  a26669a );
 a1142a <=( a26660a  and  a26649a );
 a1143a <=( a26640a  and  a26629a );
 a1144a <=( a26620a  and  a26609a );
 a1145a <=( a26600a  and  a26589a );
 a1146a <=( a26580a  and  a26569a );
 a1147a <=( a26560a  and  a26549a );
 a1148a <=( a26540a  and  a26529a );
 a1149a <=( a26520a  and  a26509a );
 a1150a <=( a26500a  and  a26489a );
 a1151a <=( a26480a  and  a26469a );
 a1152a <=( a26460a  and  a26449a );
 a1153a <=( a26440a  and  a26429a );
 a1154a <=( a26420a  and  a26409a );
 a1155a <=( a26400a  and  a26389a );
 a1156a <=( a26380a  and  a26369a );
 a1157a <=( a26360a  and  a26349a );
 a1158a <=( a26340a  and  a26329a );
 a1159a <=( a26320a  and  a26309a );
 a1160a <=( a26300a  and  a26289a );
 a1161a <=( a26280a  and  a26269a );
 a1162a <=( a26260a  and  a26249a );
 a1163a <=( a26240a  and  a26229a );
 a1164a <=( a26220a  and  a26209a );
 a1165a <=( a26200a  and  a26189a );
 a1166a <=( a26180a  and  a26169a );
 a1167a <=( a26160a  and  a26149a );
 a1168a <=( a26140a  and  a26129a );
 a1169a <=( a26120a  and  a26109a );
 a1170a <=( a26100a  and  a26089a );
 a1171a <=( a26080a  and  a26069a );
 a1172a <=( a26060a  and  a26049a );
 a1173a <=( a26040a  and  a26029a );
 a1174a <=( a26020a  and  a26009a );
 a1175a <=( a26000a  and  a25989a );
 a1176a <=( a25980a  and  a25969a );
 a1177a <=( a25960a  and  a25949a );
 a1178a <=( a25940a  and  a25929a );
 a1179a <=( a25920a  and  a25909a );
 a1180a <=( a25900a  and  a25889a );
 a1181a <=( a25880a  and  a25869a );
 a1182a <=( a25860a  and  a25849a );
 a1183a <=( a25840a  and  a25829a );
 a1184a <=( a25820a  and  a25809a );
 a1185a <=( a25800a  and  a25789a );
 a1186a <=( a25780a  and  a25769a );
 a1187a <=( a25760a  and  a25749a );
 a1188a <=( a25740a  and  a25729a );
 a1189a <=( a25720a  and  a25709a );
 a1190a <=( a25700a  and  a25689a );
 a1191a <=( a25680a  and  a25669a );
 a1192a <=( a25660a  and  a25649a );
 a1193a <=( a25640a  and  a25629a );
 a1194a <=( a25620a  and  a25609a );
 a1195a <=( a25600a  and  a25589a );
 a1196a <=( a25580a  and  a25569a );
 a1197a <=( a25560a  and  a25549a );
 a1198a <=( a25540a  and  a25529a );
 a1199a <=( a25520a  and  a25509a );
 a1200a <=( a25500a  and  a25489a );
 a1201a <=( a25480a  and  a25469a );
 a1202a <=( a25460a  and  a25449a );
 a1203a <=( a25440a  and  a25429a );
 a1204a <=( a25420a  and  a25409a );
 a1205a <=( a25400a  and  a25389a );
 a1206a <=( a25380a  and  a25369a );
 a1207a <=( a25360a  and  a25349a );
 a1208a <=( a25340a  and  a25329a );
 a1209a <=( a25320a  and  a25309a );
 a1210a <=( a25300a  and  a25289a );
 a1211a <=( a25280a  and  a25269a );
 a1212a <=( a25260a  and  a25249a );
 a1213a <=( a25240a  and  a25229a );
 a1214a <=( a25220a  and  a25209a );
 a1215a <=( a25200a  and  a25189a );
 a1216a <=( a25180a  and  a25169a );
 a1217a <=( a25160a  and  a25149a );
 a1218a <=( a25140a  and  a25129a );
 a1219a <=( a25120a  and  a25109a );
 a1220a <=( a25100a  and  a25089a );
 a1221a <=( a25080a  and  a25069a );
 a1222a <=( a25060a  and  a25049a );
 a1223a <=( a25040a  and  a25029a );
 a1224a <=( a25020a  and  a25009a );
 a1225a <=( a25000a  and  a24989a );
 a1226a <=( a24980a  and  a24969a );
 a1227a <=( a24960a  and  a24949a );
 a1228a <=( a24940a  and  a24929a );
 a1229a <=( a24920a  and  a24909a );
 a1230a <=( a24900a  and  a24889a );
 a1231a <=( a24880a  and  a24869a );
 a1232a <=( a24860a  and  a24849a );
 a1233a <=( a24840a  and  a24829a );
 a1234a <=( a24820a  and  a24809a );
 a1235a <=( a24800a  and  a24789a );
 a1236a <=( a24780a  and  a24769a );
 a1237a <=( a24760a  and  a24749a );
 a1238a <=( a24740a  and  a24729a );
 a1239a <=( a24720a  and  a24709a );
 a1240a <=( a24700a  and  a24689a );
 a1241a <=( a24680a  and  a24669a );
 a1242a <=( a24660a  and  a24649a );
 a1243a <=( a24640a  and  a24629a );
 a1244a <=( a24620a  and  a24609a );
 a1245a <=( a24600a  and  a24589a );
 a1246a <=( a24580a  and  a24569a );
 a1247a <=( a24560a  and  a24549a );
 a1248a <=( a24540a  and  a24529a );
 a1249a <=( a24520a  and  a24509a );
 a1250a <=( a24500a  and  a24489a );
 a1251a <=( a24480a  and  a24469a );
 a1252a <=( a24460a  and  a24449a );
 a1253a <=( a24440a  and  a24429a );
 a1254a <=( a24420a  and  a24409a );
 a1255a <=( a24400a  and  a24389a );
 a1256a <=( a24380a  and  a24369a );
 a1257a <=( a24360a  and  a24349a );
 a1258a <=( a24340a  and  a24329a );
 a1259a <=( a24320a  and  a24309a );
 a1260a <=( a24300a  and  a24289a );
 a1261a <=( a24280a  and  a24269a );
 a1262a <=( a24260a  and  a24249a );
 a1263a <=( a24240a  and  a24229a );
 a1264a <=( a24220a  and  a24209a );
 a1265a <=( a24200a  and  a24189a );
 a1266a <=( a24180a  and  a24169a );
 a1267a <=( a24160a  and  a24149a );
 a1268a <=( a24140a  and  a24129a );
 a1269a <=( a24120a  and  a24109a );
 a1270a <=( a24100a  and  a24089a );
 a1271a <=( a24080a  and  a24069a );
 a1272a <=( a24060a  and  a24049a );
 a1273a <=( a24040a  and  a24029a );
 a1274a <=( a24020a  and  a24009a );
 a1275a <=( a24000a  and  a23989a );
 a1276a <=( a23980a  and  a23969a );
 a1277a <=( a23960a  and  a23949a );
 a1278a <=( a23940a  and  a23929a );
 a1279a <=( a23920a  and  a23909a );
 a1280a <=( a23900a  and  a23889a );
 a1281a <=( a23880a  and  a23869a );
 a1282a <=( a23860a  and  a23849a );
 a1283a <=( a23840a  and  a23829a );
 a1284a <=( a23820a  and  a23809a );
 a1285a <=( a23800a  and  a23789a );
 a1286a <=( a23780a  and  a23769a );
 a1287a <=( a23760a  and  a23749a );
 a1288a <=( a23740a  and  a23729a );
 a1289a <=( a23720a  and  a23709a );
 a1290a <=( a23700a  and  a23689a );
 a1291a <=( a23680a  and  a23669a );
 a1292a <=( a23660a  and  a23649a );
 a1293a <=( a23640a  and  a23629a );
 a1294a <=( a23620a  and  a23609a );
 a1295a <=( a23600a  and  a23589a );
 a1296a <=( a23580a  and  a23569a );
 a1297a <=( a23560a  and  a23549a );
 a1298a <=( a23540a  and  a23529a );
 a1299a <=( a23520a  and  a23509a );
 a1300a <=( a23500a  and  a23489a );
 a1301a <=( a23480a  and  a23469a );
 a1302a <=( a23460a  and  a23449a );
 a1303a <=( a23440a  and  a23429a );
 a1304a <=( a23420a  and  a23409a );
 a1305a <=( a23400a  and  a23389a );
 a1306a <=( a23380a  and  a23369a );
 a1307a <=( a23360a  and  a23349a );
 a1308a <=( a23340a  and  a23329a );
 a1309a <=( a23320a  and  a23309a );
 a1310a <=( a23300a  and  a23289a );
 a1311a <=( a23280a  and  a23269a );
 a1312a <=( a23260a  and  a23249a );
 a1313a <=( a23240a  and  a23229a );
 a1314a <=( a23220a  and  a23209a );
 a1315a <=( a23200a  and  a23189a );
 a1316a <=( a23180a  and  a23169a );
 a1317a <=( a23160a  and  a23149a );
 a1318a <=( a23140a  and  a23129a );
 a1319a <=( a23120a  and  a23109a );
 a1320a <=( a23100a  and  a23089a );
 a1321a <=( a23080a  and  a23069a );
 a1322a <=( a23060a  and  a23049a );
 a1323a <=( a23040a  and  a23029a );
 a1324a <=( a23020a  and  a23009a );
 a1325a <=( a23000a  and  a22989a );
 a1326a <=( a22980a  and  a22969a );
 a1327a <=( a22960a  and  a22949a );
 a1328a <=( a22940a  and  a22929a );
 a1329a <=( a22920a  and  a22909a );
 a1330a <=( a22900a  and  a22889a );
 a1331a <=( a22880a  and  a22869a );
 a1332a <=( a22860a  and  a22849a );
 a1333a <=( a22840a  and  a22829a );
 a1334a <=( a22820a  and  a22809a );
 a1335a <=( a22800a  and  a22789a );
 a1336a <=( a22780a  and  a22769a );
 a1337a <=( a22760a  and  a22749a );
 a1338a <=( a22740a  and  a22729a );
 a1339a <=( a22720a  and  a22711a );
 a1340a <=( a22702a  and  a22693a );
 a1341a <=( a22684a  and  a22675a );
 a1342a <=( a22666a  and  a22657a );
 a1343a <=( a22648a  and  a22639a );
 a1344a <=( a22630a  and  a22621a );
 a1345a <=( a22612a  and  a22603a );
 a1346a <=( a22594a  and  a22585a );
 a1347a <=( a22576a  and  a22567a );
 a1348a <=( a22558a  and  a22549a );
 a1349a <=( a22540a  and  a22531a );
 a1350a <=( a22522a  and  a22513a );
 a1351a <=( a22504a  and  a22495a );
 a1352a <=( a22486a  and  a22477a );
 a1353a <=( a22468a  and  a22459a );
 a1354a <=( a22450a  and  a22441a );
 a1355a <=( a22432a  and  a22423a );
 a1356a <=( a22414a  and  a22405a );
 a1357a <=( a22396a  and  a22387a );
 a1358a <=( a22378a  and  a22369a );
 a1359a <=( a22360a  and  a22351a );
 a1360a <=( a22342a  and  a22333a );
 a1361a <=( a22324a  and  a22315a );
 a1362a <=( a22306a  and  a22297a );
 a1363a <=( a22288a  and  a22279a );
 a1364a <=( a22270a  and  a22261a );
 a1365a <=( a22252a  and  a22243a );
 a1366a <=( a22234a  and  a22225a );
 a1367a <=( a22216a  and  a22207a );
 a1368a <=( a22198a  and  a22189a );
 a1369a <=( a22180a  and  a22171a );
 a1370a <=( a22162a  and  a22153a );
 a1371a <=( a22144a  and  a22135a );
 a1372a <=( a22126a  and  a22117a );
 a1373a <=( a22108a  and  a22099a );
 a1374a <=( a22090a  and  a22081a );
 a1375a <=( a22072a  and  a22063a );
 a1376a <=( a22054a  and  a22045a );
 a1377a <=( a22036a  and  a22027a );
 a1378a <=( a22018a  and  a22009a );
 a1379a <=( a22000a  and  a21991a );
 a1380a <=( a21982a  and  a21973a );
 a1381a <=( a21964a  and  a21955a );
 a1382a <=( a21946a  and  a21937a );
 a1383a <=( a21928a  and  a21919a );
 a1384a <=( a21910a  and  a21901a );
 a1385a <=( a21892a  and  a21883a );
 a1386a <=( a21874a  and  a21865a );
 a1387a <=( a21856a  and  a21847a );
 a1388a <=( a21838a  and  a21829a );
 a1389a <=( a21820a  and  a21811a );
 a1390a <=( a21802a  and  a21793a );
 a1391a <=( a21784a  and  a21775a );
 a1392a <=( a21766a  and  a21757a );
 a1393a <=( a21748a  and  a21739a );
 a1394a <=( a21730a  and  a21721a );
 a1395a <=( a21712a  and  a21703a );
 a1396a <=( a21694a  and  a21685a );
 a1397a <=( a21676a  and  a21667a );
 a1398a <=( a21658a  and  a21649a );
 a1399a <=( a21640a  and  a21631a );
 a1400a <=( a21622a  and  a21613a );
 a1401a <=( a21604a  and  a21595a );
 a1402a <=( a21586a  and  a21577a );
 a1403a <=( a21568a  and  a21559a );
 a1404a <=( a21550a  and  a21541a );
 a1405a <=( a21532a  and  a21523a );
 a1406a <=( a21514a  and  a21505a );
 a1407a <=( a21496a  and  a21487a );
 a1408a <=( a21478a  and  a21469a );
 a1409a <=( a21460a  and  a21451a );
 a1410a <=( a21442a  and  a21433a );
 a1411a <=( a21424a  and  a21415a );
 a1412a <=( a21406a  and  a21397a );
 a1413a <=( a21388a  and  a21379a );
 a1414a <=( a21370a  and  a21361a );
 a1415a <=( a21352a  and  a21343a );
 a1416a <=( a21334a  and  a21325a );
 a1417a <=( a21316a  and  a21307a );
 a1418a <=( a21298a  and  a21289a );
 a1419a <=( a21280a  and  a21271a );
 a1420a <=( a21262a  and  a21253a );
 a1421a <=( a21244a  and  a21235a );
 a1422a <=( a21226a  and  a21217a );
 a1423a <=( a21208a  and  a21199a );
 a1424a <=( a21190a  and  a21181a );
 a1425a <=( a21172a  and  a21163a );
 a1426a <=( a21154a  and  a21145a );
 a1427a <=( a21136a  and  a21127a );
 a1428a <=( a21118a  and  a21109a );
 a1429a <=( a21100a  and  a21091a );
 a1430a <=( a21082a  and  a21073a );
 a1431a <=( a21064a  and  a21055a );
 a1432a <=( a21046a  and  a21037a );
 a1433a <=( a21028a  and  a21019a );
 a1434a <=( a21010a  and  a21001a );
 a1435a <=( a20992a  and  a20983a );
 a1436a <=( a20974a  and  a20965a );
 a1437a <=( a20956a  and  a20947a );
 a1438a <=( a20938a  and  a20929a );
 a1439a <=( a20920a  and  a20911a );
 a1440a <=( a20902a  and  a20893a );
 a1441a <=( a20884a  and  a20875a );
 a1442a <=( a20866a  and  a20857a );
 a1443a <=( a20848a  and  a20839a );
 a1444a <=( a20830a  and  a20821a );
 a1445a <=( a20812a  and  a20803a );
 a1446a <=( a20794a  and  a20785a );
 a1447a <=( a20776a  and  a20767a );
 a1448a <=( a20758a  and  a20749a );
 a1449a <=( a20740a  and  a20731a );
 a1450a <=( a20722a  and  a20713a );
 a1451a <=( a20704a  and  a20695a );
 a1452a <=( a20686a  and  a20677a );
 a1453a <=( a20668a  and  a20659a );
 a1454a <=( a20650a  and  a20641a );
 a1455a <=( a20632a  and  a20623a );
 a1456a <=( a20614a  and  a20605a );
 a1457a <=( a20596a  and  a20587a );
 a1458a <=( a20578a  and  a20569a );
 a1459a <=( a20560a  and  a20551a );
 a1460a <=( a20542a  and  a20533a );
 a1461a <=( a20524a  and  a20515a );
 a1462a <=( a20506a  and  a20497a );
 a1463a <=( a20488a  and  a20479a );
 a1464a <=( a20470a  and  a20461a );
 a1465a <=( a20452a  and  a20443a );
 a1466a <=( a20434a  and  a20425a );
 a1467a <=( a20416a  and  a20407a );
 a1468a <=( a20398a  and  a20389a );
 a1469a <=( a20380a  and  a20371a );
 a1470a <=( a20362a  and  a20353a );
 a1471a <=( a20344a  and  a20335a );
 a1472a <=( a20326a  and  a20317a );
 a1473a <=( a20308a  and  a20299a );
 a1474a <=( a20290a  and  a20281a );
 a1475a <=( a20272a  and  a20263a );
 a1476a <=( a20254a  and  a20245a );
 a1477a <=( a20236a  and  a20227a );
 a1478a <=( a20218a  and  a20209a );
 a1479a <=( a20200a  and  a20191a );
 a1480a <=( a20182a  and  a20173a );
 a1481a <=( a20164a  and  a20155a );
 a1482a <=( a20146a  and  a20137a );
 a1483a <=( a20128a  and  a20119a );
 a1484a <=( a20110a  and  a20101a );
 a1485a <=( a20092a  and  a20083a );
 a1486a <=( a20074a  and  a20065a );
 a1487a <=( a20056a  and  a20047a );
 a1488a <=( a20038a  and  a20029a );
 a1489a <=( a20020a  and  a20011a );
 a1490a <=( a20002a  and  a19993a );
 a1491a <=( a19984a  and  a19975a );
 a1492a <=( a19966a  and  a19957a );
 a1493a <=( a19948a  and  a19939a );
 a1494a <=( a19930a  and  a19921a );
 a1495a <=( a19912a  and  a19903a );
 a1496a <=( a19894a  and  a19885a );
 a1497a <=( a19876a  and  a19867a );
 a1498a <=( a19858a  and  a19849a );
 a1499a <=( a19840a  and  a19831a );
 a1500a <=( a19822a  and  a19813a );
 a1501a <=( a19804a  and  a19795a );
 a1502a <=( a19786a  and  a19777a );
 a1503a <=( a19768a  and  a19759a );
 a1504a <=( a19750a  and  a19741a );
 a1505a <=( a19732a  and  a19723a );
 a1506a <=( a19714a  and  a19705a );
 a1507a <=( a19696a  and  a19687a );
 a1508a <=( a19678a  and  a19669a );
 a1509a <=( a19660a  and  a19651a );
 a1510a <=( a19642a  and  a19633a );
 a1511a <=( a19624a  and  a19615a );
 a1512a <=( a19606a  and  a19597a );
 a1513a <=( a19588a  and  a19579a );
 a1514a <=( a19570a  and  a19561a );
 a1515a <=( a19552a  and  a19543a );
 a1516a <=( a19534a  and  a19525a );
 a1517a <=( a19516a  and  a19507a );
 a1518a <=( a19498a  and  a19489a );
 a1519a <=( a19480a  and  a19471a );
 a1520a <=( a19462a  and  a19453a );
 a1521a <=( a19444a  and  a19435a );
 a1522a <=( a19426a  and  a19417a );
 a1523a <=( a19408a  and  a19399a );
 a1524a <=( a19390a  and  a19381a );
 a1525a <=( a19372a  and  a19363a );
 a1526a <=( a19354a  and  a19345a );
 a1527a <=( a19336a  and  a19327a );
 a1528a <=( a19318a  and  a19309a );
 a1529a <=( a19300a  and  a19291a );
 a1530a <=( a19282a  and  a19273a );
 a1531a <=( a19264a  and  a19255a );
 a1532a <=( a19246a  and  a19237a );
 a1533a <=( a19228a  and  a19219a );
 a1534a <=( a19210a  and  a19201a );
 a1535a <=( a19192a  and  a19183a );
 a1536a <=( a19174a  and  a19165a );
 a1537a <=( a19156a  and  a19147a );
 a1538a <=( a19138a  and  a19129a );
 a1539a <=( a19120a  and  a19111a );
 a1540a <=( a19102a  and  a19093a );
 a1541a <=( a19084a  and  a19075a );
 a1542a <=( a19066a  and  a19057a );
 a1543a <=( a19048a  and  a19039a );
 a1544a <=( a19030a  and  a19021a );
 a1545a <=( a19012a  and  a19003a );
 a1546a <=( a18994a  and  a18985a );
 a1547a <=( a18976a  and  a18967a );
 a1548a <=( a18958a  and  a18949a );
 a1549a <=( a18940a  and  a18931a );
 a1550a <=( a18922a  and  a18913a );
 a1551a <=( a18904a  and  a18895a );
 a1552a <=( a18886a  and  a18877a );
 a1553a <=( a18868a  and  a18859a );
 a1554a <=( a18850a  and  a18841a );
 a1555a <=( a18832a  and  a18823a );
 a1556a <=( a18814a  and  a18805a );
 a1557a <=( a18796a  and  a18787a );
 a1558a <=( a18778a  and  a18769a );
 a1559a <=( a18760a  and  a18751a );
 a1560a <=( a18742a  and  a18733a );
 a1561a <=( a18724a  and  a18715a );
 a1562a <=( a18706a  and  a18697a );
 a1563a <=( a18688a  and  a18679a );
 a1564a <=( a18670a  and  a18661a );
 a1565a <=( a18652a  and  a18643a );
 a1566a <=( a18634a  and  a18625a );
 a1567a <=( a18616a  and  a18607a );
 a1568a <=( a18598a  and  a18589a );
 a1569a <=( a18580a  and  a18571a );
 a1570a <=( a18562a  and  a18553a );
 a1571a <=( a18544a  and  a18535a );
 a1572a <=( a18526a  and  a18517a );
 a1573a <=( a18508a  and  a18499a );
 a1574a <=( a18490a  and  a18481a );
 a1575a <=( a18472a  and  a18463a );
 a1576a <=( a18454a  and  a18445a );
 a1577a <=( a18436a  and  a18427a );
 a1578a <=( a18418a  and  a18409a );
 a1579a <=( a18400a  and  a18391a );
 a1580a <=( a18382a  and  a18373a );
 a1581a <=( a18364a  and  a18355a );
 a1582a <=( a18346a  and  a18337a );
 a1583a <=( a18328a  and  a18319a );
 a1584a <=( a18310a  and  a18301a );
 a1585a <=( a18292a  and  a18283a );
 a1586a <=( a18274a  and  a18265a );
 a1587a <=( a18256a  and  a18247a );
 a1588a <=( a18238a  and  a18229a );
 a1589a <=( a18220a  and  a18211a );
 a1590a <=( a18202a  and  a18193a );
 a1591a <=( a18184a  and  a18175a );
 a1592a <=( a18166a  and  a18157a );
 a1593a <=( a18148a  and  a18139a );
 a1594a <=( a18130a  and  a18121a );
 a1595a <=( a18112a  and  a18103a );
 a1596a <=( a18094a  and  a18085a );
 a1597a <=( a18076a  and  a18067a );
 a1598a <=( a18058a  and  a18049a );
 a1599a <=( a18040a  and  a18031a );
 a1600a <=( a18022a  and  a18013a );
 a1601a <=( a18004a  and  a17995a );
 a1602a <=( a17986a  and  a17977a );
 a1603a <=( a17968a  and  a17959a );
 a1604a <=( a17950a  and  a17941a );
 a1605a <=( a17932a  and  a17923a );
 a1606a <=( a17914a  and  a17905a );
 a1607a <=( a17896a  and  a17887a );
 a1608a <=( a17878a  and  a17869a );
 a1609a <=( a17860a  and  a17851a );
 a1610a <=( a17842a  and  a17833a );
 a1611a <=( a17824a  and  a17815a );
 a1612a <=( a17806a  and  a17797a );
 a1613a <=( a17788a  and  a17779a );
 a1614a <=( a17770a  and  a17761a );
 a1615a <=( a17752a  and  a17743a );
 a1616a <=( a17734a  and  a17725a );
 a1617a <=( a17716a  and  a17707a );
 a1618a <=( a17698a  and  a17689a );
 a1619a <=( a17680a  and  a17671a );
 a1620a <=( a17662a  and  a17653a );
 a1621a <=( a17644a  and  a17635a );
 a1622a <=( a17626a  and  a17617a );
 a1623a <=( a17608a  and  a17599a );
 a1624a <=( a17590a  and  a17581a );
 a1625a <=( a17572a  and  a17563a );
 a1626a <=( a17554a  and  a17545a );
 a1627a <=( a17536a  and  a17527a );
 a1628a <=( a17518a  and  a17509a );
 a1629a <=( a17500a  and  a17491a );
 a1630a <=( a17482a  and  a17473a );
 a1631a <=( a17464a  and  a17455a );
 a1632a <=( a17446a  and  a17437a );
 a1633a <=( a17428a  and  a17419a );
 a1634a <=( a17410a  and  a17401a );
 a1635a <=( a17392a  and  a17383a );
 a1636a <=( a17374a  and  a17365a );
 a1637a <=( a17356a  and  a17347a );
 a1638a <=( a17338a  and  a17329a );
 a1639a <=( a17320a  and  a17311a );
 a1640a <=( a17302a  and  a17293a );
 a1641a <=( a17284a  and  a17275a );
 a1642a <=( a17266a  and  a17257a );
 a1643a <=( a17248a  and  a17239a );
 a1644a <=( a17230a  and  a17221a );
 a1645a <=( a17212a  and  a17203a );
 a1646a <=( a17194a  and  a17185a );
 a1647a <=( a17176a  and  a17167a );
 a1648a <=( a17158a  and  a17149a );
 a1649a <=( a17140a  and  a17131a );
 a1650a <=( a17122a  and  a17113a );
 a1651a <=( a17104a  and  a17095a );
 a1652a <=( a17086a  and  a17077a );
 a1653a <=( a17068a  and  a17059a );
 a1654a <=( a17050a  and  a17041a );
 a1655a <=( a17032a  and  a17023a );
 a1656a <=( a17014a  and  a17005a );
 a1657a <=( a16996a  and  a16987a );
 a1658a <=( a16978a  and  a16969a );
 a1659a <=( a16960a  and  a16951a );
 a1660a <=( a16942a  and  a16933a );
 a1661a <=( a16924a  and  a16915a );
 a1662a <=( a16906a  and  a16897a );
 a1663a <=( a16888a  and  a16879a );
 a1664a <=( a16870a  and  a16861a );
 a1665a <=( a16852a  and  a16843a );
 a1666a <=( a16834a  and  a16825a );
 a1667a <=( a16816a  and  a16807a );
 a1668a <=( a16798a  and  a16789a );
 a1669a <=( a16780a  and  a16771a );
 a1670a <=( a16762a  and  a16753a );
 a1671a <=( a16744a  and  a16735a );
 a1672a <=( a16726a  and  a16717a );
 a1673a <=( a16708a  and  a16699a );
 a1674a <=( a16690a  and  a16681a );
 a1675a <=( a16672a  and  a16663a );
 a1676a <=( a16654a  and  a16645a );
 a1677a <=( a16636a  and  a16627a );
 a1678a <=( a16618a  and  a16609a );
 a1679a <=( a16600a  and  a16591a );
 a1680a <=( a16582a  and  a16573a );
 a1681a <=( a16564a  and  a16555a );
 a1682a <=( a16546a  and  a16537a );
 a1683a <=( a16528a  and  a16519a );
 a1684a <=( a16510a  and  a16501a );
 a1685a <=( a16492a  and  a16483a );
 a1686a <=( a16474a  and  a16465a );
 a1687a <=( a16456a  and  a16447a );
 a1688a <=( a16438a  and  a16429a );
 a1689a <=( a16420a  and  a16411a );
 a1690a <=( a16402a  and  a16393a );
 a1691a <=( a16384a  and  a16375a );
 a1692a <=( a16366a  and  a16357a );
 a1693a <=( a16348a  and  a16339a );
 a1694a <=( a16330a  and  a16321a );
 a1695a <=( a16312a  and  a16303a );
 a1696a <=( a16294a  and  a16285a );
 a1697a <=( a16276a  and  a16267a );
 a1698a <=( a16258a  and  a16249a );
 a1699a <=( a16240a  and  a16231a );
 a1700a <=( a16222a  and  a16213a );
 a1701a <=( a16204a  and  a16195a );
 a1702a <=( a16186a  and  a16177a );
 a1703a <=( a16168a  and  a16159a );
 a1704a <=( a16150a  and  a16141a );
 a1705a <=( a16132a  and  a16123a );
 a1706a <=( a16114a  and  a16105a );
 a1707a <=( a16096a  and  a16087a );
 a1708a <=( a16078a  and  a16069a );
 a1709a <=( a16060a  and  a16051a );
 a1710a <=( a16042a  and  a16033a );
 a1711a <=( a16024a  and  a16015a );
 a1712a <=( a16006a  and  a15997a );
 a1713a <=( a15988a  and  a15979a );
 a1714a <=( a15970a  and  a15961a );
 a1715a <=( a15952a  and  a15943a );
 a1716a <=( a15934a  and  a15925a );
 a1717a <=( a15916a  and  a15907a );
 a1718a <=( a15898a  and  a15889a );
 a1719a <=( a15880a  and  a15871a );
 a1720a <=( a15862a  and  a15853a );
 a1721a <=( a15844a  and  a15835a );
 a1722a <=( a15826a  and  a15817a );
 a1723a <=( a15808a  and  a15799a );
 a1724a <=( a15790a  and  a15781a );
 a1725a <=( a15772a  and  a15763a );
 a1726a <=( a15754a  and  a15745a );
 a1727a <=( a15736a  and  a15727a );
 a1728a <=( a15718a  and  a15709a );
 a1729a <=( a15700a  and  a15691a );
 a1730a <=( a15682a  and  a15673a );
 a1731a <=( a15664a  and  a15655a );
 a1732a <=( a15646a  and  a15637a );
 a1733a <=( a15628a  and  a15619a );
 a1734a <=( a15610a  and  a15601a );
 a1735a <=( a15592a  and  a15583a );
 a1736a <=( a15574a  and  a15565a );
 a1737a <=( a15556a  and  a15547a );
 a1738a <=( a15538a  and  a15529a );
 a1739a <=( a15520a  and  a15511a );
 a1740a <=( a15502a  and  a15493a );
 a1741a <=( a15484a  and  a15475a );
 a1742a <=( a15466a  and  a15457a );
 a1743a <=( a15448a  and  a15439a );
 a1744a <=( a15430a  and  a15421a );
 a1745a <=( a15412a  and  a15403a );
 a1746a <=( a15394a  and  a15385a );
 a1747a <=( a15376a  and  a15367a );
 a1748a <=( a15358a  and  a15349a );
 a1749a <=( a15340a  and  a15331a );
 a1750a <=( a15322a  and  a15313a );
 a1751a <=( a15304a  and  a15295a );
 a1752a <=( a15286a  and  a15277a );
 a1753a <=( a15268a  and  a15259a );
 a1754a <=( a15250a  and  a15241a );
 a1755a <=( a15232a  and  a15223a );
 a1756a <=( a15216a  and  a15207a );
 a1757a <=( a15200a  and  a15191a );
 a1758a <=( a15184a  and  a15175a );
 a1759a <=( a15168a  and  a15159a );
 a1760a <=( a15152a  and  a15143a );
 a1761a <=( a15136a  and  a15127a );
 a1762a <=( a15120a  and  a15111a );
 a1763a <=( a15104a  and  a15095a );
 a1764a <=( a15088a  and  a15079a );
 a1765a <=( a15072a  and  a15063a );
 a1766a <=( a15056a  and  a15047a );
 a1767a <=( a15040a  and  a15031a );
 a1768a <=( a15024a  and  a15015a );
 a1769a <=( a15008a  and  a14999a );
 a1770a <=( a14992a  and  a14983a );
 a1771a <=( a14976a  and  a14967a );
 a1772a <=( a14960a  and  a14951a );
 a1773a <=( a14944a  and  a14935a );
 a1774a <=( a14928a  and  a14919a );
 a1775a <=( a14912a  and  a14903a );
 a1776a <=( a14896a  and  a14887a );
 a1777a <=( a14880a  and  a14871a );
 a1778a <=( a14864a  and  a14855a );
 a1779a <=( a14848a  and  a14839a );
 a1780a <=( a14832a  and  a14823a );
 a1781a <=( a14816a  and  a14807a );
 a1782a <=( a14800a  and  a14791a );
 a1783a <=( a14784a  and  a14775a );
 a1784a <=( a14768a  and  a14759a );
 a1785a <=( a14752a  and  a14743a );
 a1786a <=( a14736a  and  a14727a );
 a1787a <=( a14720a  and  a14711a );
 a1788a <=( a14704a  and  a14695a );
 a1789a <=( a14688a  and  a14679a );
 a1790a <=( a14672a  and  a14663a );
 a1791a <=( a14656a  and  a14647a );
 a1792a <=( a14640a  and  a14631a );
 a1793a <=( a14624a  and  a14615a );
 a1794a <=( a14608a  and  a14599a );
 a1795a <=( a14592a  and  a14583a );
 a1796a <=( a14576a  and  a14567a );
 a1797a <=( a14560a  and  a14551a );
 a1798a <=( a14544a  and  a14535a );
 a1799a <=( a14528a  and  a14519a );
 a1800a <=( a14512a  and  a14503a );
 a1801a <=( a14496a  and  a14487a );
 a1802a <=( a14480a  and  a14471a );
 a1803a <=( a14464a  and  a14455a );
 a1804a <=( a14448a  and  a14439a );
 a1805a <=( a14432a  and  a14423a );
 a1806a <=( a14416a  and  a14407a );
 a1807a <=( a14400a  and  a14391a );
 a1808a <=( a14384a  and  a14375a );
 a1809a <=( a14368a  and  a14359a );
 a1810a <=( a14352a  and  a14343a );
 a1811a <=( a14336a  and  a14327a );
 a1812a <=( a14320a  and  a14311a );
 a1813a <=( a14304a  and  a14295a );
 a1814a <=( a14288a  and  a14279a );
 a1815a <=( a14272a  and  a14263a );
 a1816a <=( a14256a  and  a14247a );
 a1817a <=( a14240a  and  a14231a );
 a1818a <=( a14224a  and  a14215a );
 a1819a <=( a14208a  and  a14199a );
 a1820a <=( a14192a  and  a14183a );
 a1821a <=( a14176a  and  a14167a );
 a1822a <=( a14160a  and  a14151a );
 a1823a <=( a14144a  and  a14135a );
 a1824a <=( a14128a  and  a14119a );
 a1825a <=( a14112a  and  a14103a );
 a1826a <=( a14096a  and  a14087a );
 a1827a <=( a14080a  and  a14071a );
 a1828a <=( a14064a  and  a14055a );
 a1829a <=( a14048a  and  a14039a );
 a1830a <=( a14032a  and  a14023a );
 a1831a <=( a14016a  and  a14007a );
 a1832a <=( a14000a  and  a13991a );
 a1833a <=( a13984a  and  a13975a );
 a1834a <=( a13968a  and  a13959a );
 a1835a <=( a13952a  and  a13943a );
 a1836a <=( a13936a  and  a13927a );
 a1837a <=( a13920a  and  a13911a );
 a1838a <=( a13904a  and  a13895a );
 a1839a <=( a13888a  and  a13879a );
 a1840a <=( a13872a  and  a13863a );
 a1841a <=( a13856a  and  a13847a );
 a1842a <=( a13840a  and  a13831a );
 a1843a <=( a13824a  and  a13815a );
 a1844a <=( a13808a  and  a13799a );
 a1845a <=( a13792a  and  a13783a );
 a1846a <=( a13776a  and  a13767a );
 a1847a <=( a13760a  and  a13751a );
 a1848a <=( a13744a  and  a13735a );
 a1849a <=( a13728a  and  a13719a );
 a1850a <=( a13712a  and  a13703a );
 a1851a <=( a13696a  and  a13687a );
 a1852a <=( a13680a  and  a13671a );
 a1853a <=( a13664a  and  a13655a );
 a1854a <=( a13648a  and  a13639a );
 a1855a <=( a13632a  and  a13623a );
 a1856a <=( a13616a  and  a13607a );
 a1857a <=( a13600a  and  a13591a );
 a1858a <=( a13584a  and  a13575a );
 a1859a <=( a13568a  and  a13559a );
 a1860a <=( a13552a  and  a13543a );
 a1861a <=( a13536a  and  a13527a );
 a1862a <=( a13520a  and  a13511a );
 a1863a <=( a13504a  and  a13495a );
 a1864a <=( a13488a  and  a13479a );
 a1865a <=( a13472a  and  a13463a );
 a1866a <=( a13456a  and  a13447a );
 a1867a <=( a13440a  and  a13431a );
 a1868a <=( a13424a  and  a13415a );
 a1869a <=( a13408a  and  a13399a );
 a1870a <=( a13392a  and  a13383a );
 a1871a <=( a13376a  and  a13367a );
 a1872a <=( a13360a  and  a13351a );
 a1873a <=( a13344a  and  a13335a );
 a1874a <=( a13328a  and  a13319a );
 a1875a <=( a13312a  and  a13303a );
 a1876a <=( a13296a  and  a13287a );
 a1877a <=( a13280a  and  a13271a );
 a1878a <=( a13264a  and  a13255a );
 a1879a <=( a13248a  and  a13239a );
 a1880a <=( a13232a  and  a13223a );
 a1881a <=( a13216a  and  a13207a );
 a1882a <=( a13200a  and  a13191a );
 a1883a <=( a13184a  and  a13175a );
 a1884a <=( a13168a  and  a13159a );
 a1885a <=( a13152a  and  a13143a );
 a1886a <=( a13136a  and  a13127a );
 a1887a <=( a13120a  and  a13111a );
 a1888a <=( a13104a  and  a13095a );
 a1889a <=( a13088a  and  a13079a );
 a1890a <=( a13072a  and  a13063a );
 a1891a <=( a13056a  and  a13047a );
 a1892a <=( a13040a  and  a13031a );
 a1893a <=( a13024a  and  a13015a );
 a1894a <=( a13008a  and  a12999a );
 a1895a <=( a12992a  and  a12983a );
 a1896a <=( a12976a  and  a12967a );
 a1897a <=( a12960a  and  a12951a );
 a1898a <=( a12944a  and  a12935a );
 a1899a <=( a12928a  and  a12919a );
 a1900a <=( a12912a  and  a12903a );
 a1901a <=( a12896a  and  a12887a );
 a1902a <=( a12880a  and  a12871a );
 a1903a <=( a12864a  and  a12855a );
 a1904a <=( a12848a  and  a12839a );
 a1905a <=( a12832a  and  a12823a );
 a1906a <=( a12816a  and  a12807a );
 a1907a <=( a12800a  and  a12791a );
 a1908a <=( a12784a  and  a12775a );
 a1909a <=( a12768a  and  a12759a );
 a1910a <=( a12752a  and  a12743a );
 a1911a <=( a12736a  and  a12727a );
 a1912a <=( a12720a  and  a12711a );
 a1913a <=( a12704a  and  a12695a );
 a1914a <=( a12688a  and  a12679a );
 a1915a <=( a12672a  and  a12663a );
 a1916a <=( a12656a  and  a12647a );
 a1917a <=( a12640a  and  a12631a );
 a1918a <=( a12624a  and  a12615a );
 a1919a <=( a12608a  and  a12599a );
 a1920a <=( a12592a  and  a12583a );
 a1921a <=( a12576a  and  a12567a );
 a1922a <=( a12560a  and  a12551a );
 a1923a <=( a12544a  and  a12535a );
 a1924a <=( a12528a  and  a12519a );
 a1925a <=( a12512a  and  a12503a );
 a1926a <=( a12496a  and  a12487a );
 a1927a <=( a12480a  and  a12471a );
 a1928a <=( a12464a  and  a12455a );
 a1929a <=( a12448a  and  a12439a );
 a1930a <=( a12432a  and  a12423a );
 a1931a <=( a12416a  and  a12407a );
 a1932a <=( a12400a  and  a12391a );
 a1933a <=( a12384a  and  a12375a );
 a1934a <=( a12368a  and  a12359a );
 a1935a <=( a12352a  and  a12343a );
 a1936a <=( a12336a  and  a12327a );
 a1937a <=( a12320a  and  a12311a );
 a1938a <=( a12304a  and  a12295a );
 a1939a <=( a12288a  and  a12279a );
 a1940a <=( a12272a  and  a12263a );
 a1941a <=( a12256a  and  a12247a );
 a1942a <=( a12240a  and  a12231a );
 a1943a <=( a12224a  and  a12215a );
 a1944a <=( a12208a  and  a12199a );
 a1945a <=( a12192a  and  a12183a );
 a1946a <=( a12176a  and  a12167a );
 a1947a <=( a12160a  and  a12151a );
 a1948a <=( a12144a  and  a12135a );
 a1949a <=( a12128a  and  a12119a );
 a1950a <=( a12112a  and  a12103a );
 a1951a <=( a12096a  and  a12087a );
 a1952a <=( a12080a  and  a12071a );
 a1953a <=( a12064a  and  a12055a );
 a1954a <=( a12048a  and  a12039a );
 a1955a <=( a12032a  and  a12023a );
 a1956a <=( a12016a  and  a12007a );
 a1957a <=( a12000a  and  a11991a );
 a1958a <=( a11984a  and  a11975a );
 a1959a <=( a11968a  and  a11959a );
 a1960a <=( a11952a  and  a11943a );
 a1961a <=( a11936a  and  a11927a );
 a1962a <=( a11920a  and  a11911a );
 a1963a <=( a11904a  and  a11895a );
 a1964a <=( a11888a  and  a11879a );
 a1965a <=( a11872a  and  a11863a );
 a1966a <=( a11856a  and  a11847a );
 a1967a <=( a11840a  and  a11831a );
 a1968a <=( a11824a  and  a11815a );
 a1969a <=( a11808a  and  a11799a );
 a1970a <=( a11792a  and  a11783a );
 a1971a <=( a11776a  and  a11767a );
 a1972a <=( a11760a  and  a11751a );
 a1973a <=( a11744a  and  a11735a );
 a1974a <=( a11728a  and  a11719a );
 a1975a <=( a11712a  and  a11703a );
 a1976a <=( a11696a  and  a11687a );
 a1977a <=( a11680a  and  a11671a );
 a1978a <=( a11664a  and  a11655a );
 a1979a <=( a11648a  and  a11639a );
 a1980a <=( a11632a  and  a11623a );
 a1981a <=( a11616a  and  a11607a );
 a1982a <=( a11600a  and  a11591a );
 a1983a <=( a11584a  and  a11575a );
 a1984a <=( a11568a  and  a11559a );
 a1985a <=( a11552a  and  a11543a );
 a1986a <=( a11536a  and  a11527a );
 a1987a <=( a11520a  and  a11511a );
 a1988a <=( a11504a  and  a11495a );
 a1989a <=( a11488a  and  a11479a );
 a1990a <=( a11472a  and  a11463a );
 a1991a <=( a11456a  and  a11447a );
 a1992a <=( a11440a  and  a11431a );
 a1993a <=( a11424a  and  a11415a );
 a1994a <=( a11408a  and  a11399a );
 a1995a <=( a11392a  and  a11383a );
 a1996a <=( a11376a  and  a11367a );
 a1997a <=( a11360a  and  a11351a );
 a1998a <=( a11344a  and  a11335a );
 a1999a <=( a11328a  and  a11319a );
 a2000a <=( a11312a  and  a11303a );
 a2001a <=( a11296a  and  a11287a );
 a2002a <=( a11280a  and  a11271a );
 a2003a <=( a11264a  and  a11255a );
 a2004a <=( a11248a  and  a11239a );
 a2005a <=( a11232a  and  a11223a );
 a2006a <=( a11216a  and  a11207a );
 a2007a <=( a11200a  and  a11191a );
 a2008a <=( a11184a  and  a11175a );
 a2009a <=( a11168a  and  a11159a );
 a2010a <=( a11152a  and  a11143a );
 a2011a <=( a11136a  and  a11127a );
 a2012a <=( a11120a  and  a11111a );
 a2013a <=( a11104a  and  a11095a );
 a2014a <=( a11088a  and  a11079a );
 a2015a <=( a11072a  and  a11063a );
 a2016a <=( a11056a  and  a11047a );
 a2017a <=( a11040a  and  a11031a );
 a2018a <=( a11024a  and  a11015a );
 a2019a <=( a11008a  and  a10999a );
 a2020a <=( a10992a  and  a10983a );
 a2021a <=( a10976a  and  a10967a );
 a2022a <=( a10960a  and  a10951a );
 a2023a <=( a10944a  and  a10935a );
 a2024a <=( a10928a  and  a10919a );
 a2025a <=( a10912a  and  a10903a );
 a2026a <=( a10896a  and  a10887a );
 a2027a <=( a10880a  and  a10871a );
 a2028a <=( a10864a  and  a10855a );
 a2029a <=( a10848a  and  a10839a );
 a2030a <=( a10832a  and  a10823a );
 a2031a <=( a10816a  and  a10807a );
 a2032a <=( a10800a  and  a10791a );
 a2033a <=( a10784a  and  a10775a );
 a2034a <=( a10768a  and  a10759a );
 a2035a <=( a10752a  and  a10743a );
 a2036a <=( a10736a  and  a10727a );
 a2037a <=( a10720a  and  a10711a );
 a2038a <=( a10704a  and  a10695a );
 a2039a <=( a10688a  and  a10679a );
 a2040a <=( a10672a  and  a10663a );
 a2041a <=( a10656a  and  a10647a );
 a2042a <=( a10640a  and  a10631a );
 a2043a <=( a10624a  and  a10615a );
 a2044a <=( a10608a  and  a10599a );
 a2045a <=( a10592a  and  a10583a );
 a2046a <=( a10576a  and  a10567a );
 a2047a <=( a10560a  and  a10551a );
 a2048a <=( a10544a  and  a10535a );
 a2049a <=( a10528a  and  a10519a );
 a2050a <=( a10512a  and  a10503a );
 a2051a <=( a10496a  and  a10487a );
 a2052a <=( a10480a  and  a10471a );
 a2053a <=( a10464a  and  a10455a );
 a2054a <=( a10448a  and  a10439a );
 a2055a <=( a10432a  and  a10423a );
 a2056a <=( a10416a  and  a10407a );
 a2057a <=( a10400a  and  a10391a );
 a2058a <=( a10384a  and  a10375a );
 a2059a <=( a10368a  and  a10359a );
 a2060a <=( a10352a  and  a10343a );
 a2061a <=( a10336a  and  a10327a );
 a2062a <=( a10320a  and  a10311a );
 a2063a <=( a10304a  and  a10295a );
 a2064a <=( a10288a  and  a10279a );
 a2065a <=( a10272a  and  a10263a );
 a2066a <=( a10256a  and  a10247a );
 a2067a <=( a10240a  and  a10231a );
 a2068a <=( a10224a  and  a10215a );
 a2069a <=( a10208a  and  a10199a );
 a2070a <=( a10192a  and  a10183a );
 a2071a <=( a10176a  and  a10167a );
 a2072a <=( a10160a  and  a10151a );
 a2073a <=( a10144a  and  a10135a );
 a2074a <=( a10128a  and  a10119a );
 a2075a <=( a10112a  and  a10103a );
 a2076a <=( a10096a  and  a10087a );
 a2077a <=( a10080a  and  a10071a );
 a2078a <=( a10064a  and  a10055a );
 a2079a <=( a10048a  and  a10039a );
 a2080a <=( a10032a  and  a10023a );
 a2081a <=( a10016a  and  a10007a );
 a2082a <=( a10000a  and  a9991a );
 a2083a <=( a9984a  and  a9977a );
 a2084a <=( a9970a  and  a9963a );
 a2085a <=( a9956a  and  a9949a );
 a2086a <=( a9942a  and  a9935a );
 a2087a <=( a9928a  and  a9921a );
 a2088a <=( a9914a  and  a9907a );
 a2089a <=( a9900a  and  a9893a );
 a2090a <=( a9886a  and  a9879a );
 a2091a <=( a9872a  and  a9865a );
 a2092a <=( a9858a  and  a9851a );
 a2093a <=( a9844a  and  a9837a );
 a2094a <=( a9830a  and  a9823a );
 a2095a <=( a9816a  and  a9809a );
 a2096a <=( a9802a  and  a9795a );
 a2097a <=( a9788a  and  a9781a );
 a2098a <=( a9774a  and  a9767a );
 a2099a <=( a9760a  and  a9753a );
 a2100a <=( a9746a  and  a9739a );
 a2101a <=( a9732a  and  a9725a );
 a2102a <=( a9718a  and  a9711a );
 a2103a <=( a9704a  and  a9697a );
 a2104a <=( a9690a  and  a9683a );
 a2105a <=( a9676a  and  a9669a );
 a2106a <=( a9662a  and  a9655a );
 a2107a <=( a9648a  and  a9641a );
 a2108a <=( a9634a  and  a9627a );
 a2109a <=( a9620a  and  a9613a );
 a2110a <=( a9606a  and  a9599a );
 a2111a <=( a9592a  and  a9585a );
 a2112a <=( a9578a  and  a9571a );
 a2113a <=( a9564a  and  a9557a );
 a2114a <=( a9550a  and  a9543a );
 a2115a <=( a9536a  and  a9529a );
 a2116a <=( a9522a  and  a9515a );
 a2117a <=( a9508a  and  a9501a );
 a2118a <=( a9494a  and  a9487a );
 a2119a <=( a9480a  and  a9473a );
 a2120a <=( a9466a  and  a9459a );
 a2121a <=( a9452a  and  a9445a );
 a2122a <=( a9438a  and  a9431a );
 a2123a <=( a9424a  and  a9417a );
 a2124a <=( a9410a  and  a9403a );
 a2125a <=( a9396a  and  a9389a );
 a2126a <=( a9382a  and  a9375a );
 a2127a <=( a9368a  and  a9361a );
 a2128a <=( a9354a  and  a9347a );
 a2129a <=( a9340a  and  a9333a );
 a2130a <=( a9326a  and  a9319a );
 a2131a <=( a9312a  and  a9305a );
 a2132a <=( a9298a  and  a9291a );
 a2133a <=( a9284a  and  a9277a );
 a2134a <=( a9270a  and  a9263a );
 a2135a <=( a9256a  and  a9249a );
 a2136a <=( a9242a  and  a9235a );
 a2137a <=( a9228a  and  a9221a );
 a2138a <=( a9214a  and  a9207a );
 a2139a <=( a9200a  and  a9193a );
 a2140a <=( a9186a  and  a9179a );
 a2141a <=( a9172a  and  a9165a );
 a2142a <=( a9158a  and  a9151a );
 a2143a <=( a9144a  and  a9137a );
 a2144a <=( a9130a  and  a9123a );
 a2145a <=( a9116a  and  a9109a );
 a2146a <=( a9102a  and  a9095a );
 a2147a <=( a9088a  and  a9081a );
 a2148a <=( a9074a  and  a9067a );
 a2149a <=( a9060a  and  a9053a );
 a2150a <=( a9046a  and  a9039a );
 a2151a <=( a9032a  and  a9025a );
 a2152a <=( a9018a  and  a9011a );
 a2153a <=( a9004a  and  a8997a );
 a2154a <=( a8990a  and  a8983a );
 a2155a <=( a8976a  and  a8969a );
 a2156a <=( a8962a  and  a8955a );
 a2157a <=( a8948a  and  a8941a );
 a2158a <=( a8934a  and  a8927a );
 a2159a <=( a8920a  and  a8913a );
 a2160a <=( a8906a  and  a8899a );
 a2161a <=( a8892a  and  a8885a );
 a2162a <=( a8878a  and  a8871a );
 a2163a <=( a8864a  and  a8857a );
 a2164a <=( a8850a  and  a8843a );
 a2165a <=( a8836a  and  a8829a );
 a2166a <=( a8822a  and  a8815a );
 a2167a <=( a8808a  and  a8801a );
 a2168a <=( a8794a  and  a8787a );
 a2169a <=( a8780a  and  a8773a );
 a2170a <=( a8766a  and  a8759a );
 a2171a <=( a8752a  and  a8745a );
 a2172a <=( a8738a  and  a8731a );
 a2173a <=( a8724a  and  a8717a );
 a2174a <=( a8710a  and  a8703a );
 a2175a <=( a8696a  and  a8689a );
 a2176a <=( a8682a  and  a8675a );
 a2177a <=( a8668a  and  a8661a );
 a2178a <=( a8654a  and  a8647a );
 a2179a <=( a8640a  and  a8633a );
 a2180a <=( a8626a  and  a8619a );
 a2181a <=( a8612a  and  a8605a );
 a2182a <=( a8598a  and  a8591a );
 a2183a <=( a8584a  and  a8577a );
 a2184a <=( a8570a  and  a8563a );
 a2185a <=( a8556a  and  a8549a );
 a2186a <=( a8542a  and  a8535a );
 a2187a <=( a8528a  and  a8521a );
 a2188a <=( a8514a  and  a8507a );
 a2189a <=( a8500a  and  a8493a );
 a2190a <=( a8486a  and  a8479a );
 a2191a <=( a8472a  and  a8465a );
 a2192a <=( a8458a  and  a8451a );
 a2193a <=( a8444a  and  a8437a );
 a2194a <=( a8430a  and  a8423a );
 a2195a <=( a8416a  and  a8409a );
 a2196a <=( a8402a  and  a8395a );
 a2197a <=( a8388a  and  a8381a );
 a2198a <=( a8374a  and  a8367a );
 a2199a <=( a8360a  and  a8353a );
 a2200a <=( a8346a  and  a8339a );
 a2201a <=( a8332a  and  a8325a );
 a2202a <=( a8318a  and  a8311a );
 a2203a <=( a8304a  and  a8297a );
 a2204a <=( a8290a  and  a8283a );
 a2205a <=( a8276a  and  a8269a );
 a2206a <=( a8262a  and  a8255a );
 a2207a <=( a8248a  and  a8241a );
 a2208a <=( a8234a  and  a8227a );
 a2209a <=( a8220a  and  a8213a );
 a2210a <=( a8206a  and  a8199a );
 a2211a <=( a8192a  and  a8185a );
 a2212a <=( a8178a  and  a8171a );
 a2213a <=( a8164a  and  a8157a );
 a2214a <=( a8150a  and  a8143a );
 a2215a <=( a8136a  and  a8129a );
 a2216a <=( a8122a  and  a8115a );
 a2217a <=( a8108a  and  a8101a );
 a2218a <=( a8094a  and  a8087a );
 a2219a <=( a8080a  and  a8073a );
 a2220a <=( a8066a  and  a8059a );
 a2221a <=( a8052a  and  a8045a );
 a2222a <=( a8038a  and  a8031a );
 a2223a <=( a8024a  and  a8017a );
 a2224a <=( a8010a  and  a8003a );
 a2225a <=( a7996a  and  a7989a );
 a2226a <=( a7982a  and  a7975a );
 a2227a <=( a7968a  and  a7961a );
 a2228a <=( a7954a  and  a7947a );
 a2229a <=( a7940a  and  a7933a );
 a2230a <=( a7926a  and  a7919a );
 a2231a <=( a7912a  and  a7905a );
 a2232a <=( a7898a  and  a7891a );
 a2233a <=( a7884a  and  a7877a );
 a2234a <=( a7870a  and  a7863a );
 a2235a <=( a7856a  and  a7849a );
 a2236a <=( a7842a  and  a7835a );
 a2237a <=( a7828a  and  a7821a );
 a2238a <=( a7814a  and  a7807a );
 a2239a <=( a7800a  and  a7793a );
 a2240a <=( a7786a  and  a7779a );
 a2241a <=( a7772a  and  a7765a );
 a2242a <=( a7758a  and  a7751a );
 a2243a <=( a7744a  and  a7737a );
 a2244a <=( a7730a  and  a7723a );
 a2245a <=( a7716a  and  a7709a );
 a2246a <=( a7702a  and  a7695a );
 a2247a <=( a7688a  and  a7681a );
 a2248a <=( a7674a  and  a7667a );
 a2249a <=( a7660a  and  a7653a );
 a2250a <=( a7646a  and  a7639a );
 a2251a <=( a7632a  and  a7625a );
 a2252a <=( a7620a  and  a7613a );
 a2253a <=( a7608a  and  a7601a );
 a2254a <=( a7596a  and  a7589a );
 a2255a <=( a7584a  and  a7577a );
 a2256a <=( a7572a  and  a7565a );
 a2257a <=( a7560a  and  a7553a );
 a2258a <=( a7548a  and  a7541a );
 a2259a <=( a7536a  and  a7529a );
 a2260a <=( a7524a  and  a7517a );
 a2261a <=( a7512a  and  a7505a );
 a2262a <=( a7500a  and  a7493a );
 a2263a <=( a7488a  and  a7481a );
 a2264a <=( a7476a  and  a7469a );
 a2265a <=( a7464a  and  a7457a );
 a2266a <=( a7452a  and  a7445a );
 a2267a <=( a7440a  and  a7433a );
 a2268a <=( a7428a  and  a7421a );
 a2269a <=( a7416a  and  a7409a );
 a2270a <=( a7404a  and  a7397a );
 a2271a <=( a7392a  and  a7385a );
 a2272a <=( a7380a  and  a7373a );
 a2273a <=( a7368a  and  a7361a );
 a2274a <=( a7356a  and  a7349a );
 a2275a <=( a7344a  and  a7337a );
 a2276a <=( a7332a  and  a7325a );
 a2277a <=( a7320a  and  a7313a );
 a2278a <=( a7308a  and  a7301a );
 a2279a <=( a7296a  and  a7289a );
 a2280a <=( a7284a  and  a7277a );
 a2281a <=( a7272a  and  a7265a );
 a2282a <=( a7260a  and  a7253a );
 a2283a <=( a7248a  and  a7241a );
 a2284a <=( a7236a  and  a7229a );
 a2285a <=( a7224a  and  a7217a );
 a2286a <=( a7212a  and  a7205a );
 a2287a <=( a7200a  and  a7193a );
 a2288a <=( a7188a  and  a7181a );
 a2289a <=( a7176a  and  a7169a );
 a2290a <=( a7164a  and  a7157a );
 a2291a <=( a7152a  and  a7145a );
 a2292a <=( a7140a  and  a7133a );
 a2293a <=( a7128a  and  a7121a );
 a2294a <=( a7116a  and  a7109a );
 a2295a <=( a7104a  and  a7097a );
 a2296a <=( a7092a  and  a7085a );
 a2297a <=( a7080a  and  a7073a );
 a2298a <=( a7068a  and  a7061a );
 a2299a <=( a7056a  and  a7049a );
 a2300a <=( a7044a  and  a7037a );
 a2301a <=( a7032a  and  a7025a );
 a2302a <=( a7020a  and  a7013a );
 a2303a <=( a7008a  and  a7003a );
 a2304a <=( a6998a  and  a6993a );
 a2305a <=( a6988a  and  a6983a );
 a2306a <=( a6978a  and  a6973a );
 a2307a <=( a6968a  and  a6963a );
 a2308a <=( a6958a  and  a6953a );
 a2309a <=( a6948a  and  a6943a );
 a2310a <=( a6938a  and  a6933a );
 a2313a <=( a2309a ) or ( a2310a );
 a2316a <=( a2307a ) or ( a2308a );
 a2317a <=( a2316a ) or ( a2313a );
 a2320a <=( a2305a ) or ( a2306a );
 a2324a <=( a2302a ) or ( a2303a );
 a2325a <=( a2304a ) or ( a2324a );
 a2326a <=( a2325a ) or ( a2320a );
 a2327a <=( a2326a ) or ( a2317a );
 a2330a <=( a2300a ) or ( a2301a );
 a2333a <=( a2298a ) or ( a2299a );
 a2334a <=( a2333a ) or ( a2330a );
 a2337a <=( a2296a ) or ( a2297a );
 a2341a <=( a2293a ) or ( a2294a );
 a2342a <=( a2295a ) or ( a2341a );
 a2343a <=( a2342a ) or ( a2337a );
 a2344a <=( a2343a ) or ( a2334a );
 a2345a <=( a2344a ) or ( a2327a );
 a2348a <=( a2291a ) or ( a2292a );
 a2351a <=( a2289a ) or ( a2290a );
 a2352a <=( a2351a ) or ( a2348a );
 a2355a <=( a2287a ) or ( a2288a );
 a2359a <=( a2284a ) or ( a2285a );
 a2360a <=( a2286a ) or ( a2359a );
 a2361a <=( a2360a ) or ( a2355a );
 a2362a <=( a2361a ) or ( a2352a );
 a2365a <=( a2282a ) or ( a2283a );
 a2368a <=( a2280a ) or ( a2281a );
 a2369a <=( a2368a ) or ( a2365a );
 a2372a <=( a2278a ) or ( a2279a );
 a2376a <=( a2275a ) or ( a2276a );
 a2377a <=( a2277a ) or ( a2376a );
 a2378a <=( a2377a ) or ( a2372a );
 a2379a <=( a2378a ) or ( a2369a );
 a2380a <=( a2379a ) or ( a2362a );
 a2381a <=( a2380a ) or ( a2345a );
 a2384a <=( a2273a ) or ( a2274a );
 a2387a <=( a2271a ) or ( a2272a );
 a2388a <=( a2387a ) or ( a2384a );
 a2391a <=( a2269a ) or ( a2270a );
 a2395a <=( a2266a ) or ( a2267a );
 a2396a <=( a2268a ) or ( a2395a );
 a2397a <=( a2396a ) or ( a2391a );
 a2398a <=( a2397a ) or ( a2388a );
 a2401a <=( a2264a ) or ( a2265a );
 a2404a <=( a2262a ) or ( a2263a );
 a2405a <=( a2404a ) or ( a2401a );
 a2408a <=( a2260a ) or ( a2261a );
 a2412a <=( a2257a ) or ( a2258a );
 a2413a <=( a2259a ) or ( a2412a );
 a2414a <=( a2413a ) or ( a2408a );
 a2415a <=( a2414a ) or ( a2405a );
 a2416a <=( a2415a ) or ( a2398a );
 a2419a <=( a2255a ) or ( a2256a );
 a2422a <=( a2253a ) or ( a2254a );
 a2423a <=( a2422a ) or ( a2419a );
 a2426a <=( a2251a ) or ( a2252a );
 a2430a <=( a2248a ) or ( a2249a );
 a2431a <=( a2250a ) or ( a2430a );
 a2432a <=( a2431a ) or ( a2426a );
 a2433a <=( a2432a ) or ( a2423a );
 a2436a <=( a2246a ) or ( a2247a );
 a2439a <=( a2244a ) or ( a2245a );
 a2440a <=( a2439a ) or ( a2436a );
 a2443a <=( a2242a ) or ( a2243a );
 a2447a <=( a2239a ) or ( a2240a );
 a2448a <=( a2241a ) or ( a2447a );
 a2449a <=( a2448a ) or ( a2443a );
 a2450a <=( a2449a ) or ( a2440a );
 a2451a <=( a2450a ) or ( a2433a );
 a2452a <=( a2451a ) or ( a2416a );
 a2453a <=( a2452a ) or ( a2381a );
 a2456a <=( a2237a ) or ( a2238a );
 a2459a <=( a2235a ) or ( a2236a );
 a2460a <=( a2459a ) or ( a2456a );
 a2463a <=( a2233a ) or ( a2234a );
 a2467a <=( a2230a ) or ( a2231a );
 a2468a <=( a2232a ) or ( a2467a );
 a2469a <=( a2468a ) or ( a2463a );
 a2470a <=( a2469a ) or ( a2460a );
 a2473a <=( a2228a ) or ( a2229a );
 a2476a <=( a2226a ) or ( a2227a );
 a2477a <=( a2476a ) or ( a2473a );
 a2480a <=( a2224a ) or ( a2225a );
 a2484a <=( a2221a ) or ( a2222a );
 a2485a <=( a2223a ) or ( a2484a );
 a2486a <=( a2485a ) or ( a2480a );
 a2487a <=( a2486a ) or ( a2477a );
 a2488a <=( a2487a ) or ( a2470a );
 a2491a <=( a2219a ) or ( a2220a );
 a2494a <=( a2217a ) or ( a2218a );
 a2495a <=( a2494a ) or ( a2491a );
 a2498a <=( a2215a ) or ( a2216a );
 a2502a <=( a2212a ) or ( a2213a );
 a2503a <=( a2214a ) or ( a2502a );
 a2504a <=( a2503a ) or ( a2498a );
 a2505a <=( a2504a ) or ( a2495a );
 a2508a <=( a2210a ) or ( a2211a );
 a2511a <=( a2208a ) or ( a2209a );
 a2512a <=( a2511a ) or ( a2508a );
 a2515a <=( a2206a ) or ( a2207a );
 a2519a <=( a2203a ) or ( a2204a );
 a2520a <=( a2205a ) or ( a2519a );
 a2521a <=( a2520a ) or ( a2515a );
 a2522a <=( a2521a ) or ( a2512a );
 a2523a <=( a2522a ) or ( a2505a );
 a2524a <=( a2523a ) or ( a2488a );
 a2527a <=( a2201a ) or ( a2202a );
 a2530a <=( a2199a ) or ( a2200a );
 a2531a <=( a2530a ) or ( a2527a );
 a2534a <=( a2197a ) or ( a2198a );
 a2538a <=( a2194a ) or ( a2195a );
 a2539a <=( a2196a ) or ( a2538a );
 a2540a <=( a2539a ) or ( a2534a );
 a2541a <=( a2540a ) or ( a2531a );
 a2544a <=( a2192a ) or ( a2193a );
 a2547a <=( a2190a ) or ( a2191a );
 a2548a <=( a2547a ) or ( a2544a );
 a2551a <=( a2188a ) or ( a2189a );
 a2555a <=( a2185a ) or ( a2186a );
 a2556a <=( a2187a ) or ( a2555a );
 a2557a <=( a2556a ) or ( a2551a );
 a2558a <=( a2557a ) or ( a2548a );
 a2559a <=( a2558a ) or ( a2541a );
 a2562a <=( a2183a ) or ( a2184a );
 a2565a <=( a2181a ) or ( a2182a );
 a2566a <=( a2565a ) or ( a2562a );
 a2569a <=( a2179a ) or ( a2180a );
 a2573a <=( a2176a ) or ( a2177a );
 a2574a <=( a2178a ) or ( a2573a );
 a2575a <=( a2574a ) or ( a2569a );
 a2576a <=( a2575a ) or ( a2566a );
 a2579a <=( a2174a ) or ( a2175a );
 a2582a <=( a2172a ) or ( a2173a );
 a2583a <=( a2582a ) or ( a2579a );
 a2586a <=( a2170a ) or ( a2171a );
 a2590a <=( a2167a ) or ( a2168a );
 a2591a <=( a2169a ) or ( a2590a );
 a2592a <=( a2591a ) or ( a2586a );
 a2593a <=( a2592a ) or ( a2583a );
 a2594a <=( a2593a ) or ( a2576a );
 a2595a <=( a2594a ) or ( a2559a );
 a2596a <=( a2595a ) or ( a2524a );
 a2597a <=( a2596a ) or ( a2453a );
 a2600a <=( a2165a ) or ( a2166a );
 a2603a <=( a2163a ) or ( a2164a );
 a2604a <=( a2603a ) or ( a2600a );
 a2607a <=( a2161a ) or ( a2162a );
 a2611a <=( a2158a ) or ( a2159a );
 a2612a <=( a2160a ) or ( a2611a );
 a2613a <=( a2612a ) or ( a2607a );
 a2614a <=( a2613a ) or ( a2604a );
 a2617a <=( a2156a ) or ( a2157a );
 a2620a <=( a2154a ) or ( a2155a );
 a2621a <=( a2620a ) or ( a2617a );
 a2624a <=( a2152a ) or ( a2153a );
 a2628a <=( a2149a ) or ( a2150a );
 a2629a <=( a2151a ) or ( a2628a );
 a2630a <=( a2629a ) or ( a2624a );
 a2631a <=( a2630a ) or ( a2621a );
 a2632a <=( a2631a ) or ( a2614a );
 a2635a <=( a2147a ) or ( a2148a );
 a2638a <=( a2145a ) or ( a2146a );
 a2639a <=( a2638a ) or ( a2635a );
 a2642a <=( a2143a ) or ( a2144a );
 a2646a <=( a2140a ) or ( a2141a );
 a2647a <=( a2142a ) or ( a2646a );
 a2648a <=( a2647a ) or ( a2642a );
 a2649a <=( a2648a ) or ( a2639a );
 a2652a <=( a2138a ) or ( a2139a );
 a2655a <=( a2136a ) or ( a2137a );
 a2656a <=( a2655a ) or ( a2652a );
 a2659a <=( a2134a ) or ( a2135a );
 a2663a <=( a2131a ) or ( a2132a );
 a2664a <=( a2133a ) or ( a2663a );
 a2665a <=( a2664a ) or ( a2659a );
 a2666a <=( a2665a ) or ( a2656a );
 a2667a <=( a2666a ) or ( a2649a );
 a2668a <=( a2667a ) or ( a2632a );
 a2671a <=( a2129a ) or ( a2130a );
 a2674a <=( a2127a ) or ( a2128a );
 a2675a <=( a2674a ) or ( a2671a );
 a2678a <=( a2125a ) or ( a2126a );
 a2682a <=( a2122a ) or ( a2123a );
 a2683a <=( a2124a ) or ( a2682a );
 a2684a <=( a2683a ) or ( a2678a );
 a2685a <=( a2684a ) or ( a2675a );
 a2688a <=( a2120a ) or ( a2121a );
 a2691a <=( a2118a ) or ( a2119a );
 a2692a <=( a2691a ) or ( a2688a );
 a2695a <=( a2116a ) or ( a2117a );
 a2699a <=( a2113a ) or ( a2114a );
 a2700a <=( a2115a ) or ( a2699a );
 a2701a <=( a2700a ) or ( a2695a );
 a2702a <=( a2701a ) or ( a2692a );
 a2703a <=( a2702a ) or ( a2685a );
 a2706a <=( a2111a ) or ( a2112a );
 a2709a <=( a2109a ) or ( a2110a );
 a2710a <=( a2709a ) or ( a2706a );
 a2713a <=( a2107a ) or ( a2108a );
 a2717a <=( a2104a ) or ( a2105a );
 a2718a <=( a2106a ) or ( a2717a );
 a2719a <=( a2718a ) or ( a2713a );
 a2720a <=( a2719a ) or ( a2710a );
 a2723a <=( a2102a ) or ( a2103a );
 a2726a <=( a2100a ) or ( a2101a );
 a2727a <=( a2726a ) or ( a2723a );
 a2730a <=( a2098a ) or ( a2099a );
 a2734a <=( a2095a ) or ( a2096a );
 a2735a <=( a2097a ) or ( a2734a );
 a2736a <=( a2735a ) or ( a2730a );
 a2737a <=( a2736a ) or ( a2727a );
 a2738a <=( a2737a ) or ( a2720a );
 a2739a <=( a2738a ) or ( a2703a );
 a2740a <=( a2739a ) or ( a2668a );
 a2743a <=( a2093a ) or ( a2094a );
 a2746a <=( a2091a ) or ( a2092a );
 a2747a <=( a2746a ) or ( a2743a );
 a2750a <=( a2089a ) or ( a2090a );
 a2754a <=( a2086a ) or ( a2087a );
 a2755a <=( a2088a ) or ( a2754a );
 a2756a <=( a2755a ) or ( a2750a );
 a2757a <=( a2756a ) or ( a2747a );
 a2760a <=( a2084a ) or ( a2085a );
 a2763a <=( a2082a ) or ( a2083a );
 a2764a <=( a2763a ) or ( a2760a );
 a2767a <=( a2080a ) or ( a2081a );
 a2771a <=( a2077a ) or ( a2078a );
 a2772a <=( a2079a ) or ( a2771a );
 a2773a <=( a2772a ) or ( a2767a );
 a2774a <=( a2773a ) or ( a2764a );
 a2775a <=( a2774a ) or ( a2757a );
 a2778a <=( a2075a ) or ( a2076a );
 a2781a <=( a2073a ) or ( a2074a );
 a2782a <=( a2781a ) or ( a2778a );
 a2785a <=( a2071a ) or ( a2072a );
 a2789a <=( a2068a ) or ( a2069a );
 a2790a <=( a2070a ) or ( a2789a );
 a2791a <=( a2790a ) or ( a2785a );
 a2792a <=( a2791a ) or ( a2782a );
 a2795a <=( a2066a ) or ( a2067a );
 a2798a <=( a2064a ) or ( a2065a );
 a2799a <=( a2798a ) or ( a2795a );
 a2802a <=( a2062a ) or ( a2063a );
 a2806a <=( a2059a ) or ( a2060a );
 a2807a <=( a2061a ) or ( a2806a );
 a2808a <=( a2807a ) or ( a2802a );
 a2809a <=( a2808a ) or ( a2799a );
 a2810a <=( a2809a ) or ( a2792a );
 a2811a <=( a2810a ) or ( a2775a );
 a2814a <=( a2057a ) or ( a2058a );
 a2817a <=( a2055a ) or ( a2056a );
 a2818a <=( a2817a ) or ( a2814a );
 a2821a <=( a2053a ) or ( a2054a );
 a2825a <=( a2050a ) or ( a2051a );
 a2826a <=( a2052a ) or ( a2825a );
 a2827a <=( a2826a ) or ( a2821a );
 a2828a <=( a2827a ) or ( a2818a );
 a2831a <=( a2048a ) or ( a2049a );
 a2834a <=( a2046a ) or ( a2047a );
 a2835a <=( a2834a ) or ( a2831a );
 a2838a <=( a2044a ) or ( a2045a );
 a2842a <=( a2041a ) or ( a2042a );
 a2843a <=( a2043a ) or ( a2842a );
 a2844a <=( a2843a ) or ( a2838a );
 a2845a <=( a2844a ) or ( a2835a );
 a2846a <=( a2845a ) or ( a2828a );
 a2849a <=( a2039a ) or ( a2040a );
 a2852a <=( a2037a ) or ( a2038a );
 a2853a <=( a2852a ) or ( a2849a );
 a2856a <=( a2035a ) or ( a2036a );
 a2860a <=( a2032a ) or ( a2033a );
 a2861a <=( a2034a ) or ( a2860a );
 a2862a <=( a2861a ) or ( a2856a );
 a2863a <=( a2862a ) or ( a2853a );
 a2866a <=( a2030a ) or ( a2031a );
 a2869a <=( a2028a ) or ( a2029a );
 a2870a <=( a2869a ) or ( a2866a );
 a2873a <=( a2026a ) or ( a2027a );
 a2877a <=( a2023a ) or ( a2024a );
 a2878a <=( a2025a ) or ( a2877a );
 a2879a <=( a2878a ) or ( a2873a );
 a2880a <=( a2879a ) or ( a2870a );
 a2881a <=( a2880a ) or ( a2863a );
 a2882a <=( a2881a ) or ( a2846a );
 a2883a <=( a2882a ) or ( a2811a );
 a2884a <=( a2883a ) or ( a2740a );
 a2885a <=( a2884a ) or ( a2597a );
 a2888a <=( a2021a ) or ( a2022a );
 a2891a <=( a2019a ) or ( a2020a );
 a2892a <=( a2891a ) or ( a2888a );
 a2895a <=( a2017a ) or ( a2018a );
 a2899a <=( a2014a ) or ( a2015a );
 a2900a <=( a2016a ) or ( a2899a );
 a2901a <=( a2900a ) or ( a2895a );
 a2902a <=( a2901a ) or ( a2892a );
 a2905a <=( a2012a ) or ( a2013a );
 a2908a <=( a2010a ) or ( a2011a );
 a2909a <=( a2908a ) or ( a2905a );
 a2912a <=( a2008a ) or ( a2009a );
 a2916a <=( a2005a ) or ( a2006a );
 a2917a <=( a2007a ) or ( a2916a );
 a2918a <=( a2917a ) or ( a2912a );
 a2919a <=( a2918a ) or ( a2909a );
 a2920a <=( a2919a ) or ( a2902a );
 a2923a <=( a2003a ) or ( a2004a );
 a2926a <=( a2001a ) or ( a2002a );
 a2927a <=( a2926a ) or ( a2923a );
 a2930a <=( a1999a ) or ( a2000a );
 a2934a <=( a1996a ) or ( a1997a );
 a2935a <=( a1998a ) or ( a2934a );
 a2936a <=( a2935a ) or ( a2930a );
 a2937a <=( a2936a ) or ( a2927a );
 a2940a <=( a1994a ) or ( a1995a );
 a2943a <=( a1992a ) or ( a1993a );
 a2944a <=( a2943a ) or ( a2940a );
 a2947a <=( a1990a ) or ( a1991a );
 a2951a <=( a1987a ) or ( a1988a );
 a2952a <=( a1989a ) or ( a2951a );
 a2953a <=( a2952a ) or ( a2947a );
 a2954a <=( a2953a ) or ( a2944a );
 a2955a <=( a2954a ) or ( a2937a );
 a2956a <=( a2955a ) or ( a2920a );
 a2959a <=( a1985a ) or ( a1986a );
 a2962a <=( a1983a ) or ( a1984a );
 a2963a <=( a2962a ) or ( a2959a );
 a2966a <=( a1981a ) or ( a1982a );
 a2970a <=( a1978a ) or ( a1979a );
 a2971a <=( a1980a ) or ( a2970a );
 a2972a <=( a2971a ) or ( a2966a );
 a2973a <=( a2972a ) or ( a2963a );
 a2976a <=( a1976a ) or ( a1977a );
 a2979a <=( a1974a ) or ( a1975a );
 a2980a <=( a2979a ) or ( a2976a );
 a2983a <=( a1972a ) or ( a1973a );
 a2987a <=( a1969a ) or ( a1970a );
 a2988a <=( a1971a ) or ( a2987a );
 a2989a <=( a2988a ) or ( a2983a );
 a2990a <=( a2989a ) or ( a2980a );
 a2991a <=( a2990a ) or ( a2973a );
 a2994a <=( a1967a ) or ( a1968a );
 a2997a <=( a1965a ) or ( a1966a );
 a2998a <=( a2997a ) or ( a2994a );
 a3001a <=( a1963a ) or ( a1964a );
 a3005a <=( a1960a ) or ( a1961a );
 a3006a <=( a1962a ) or ( a3005a );
 a3007a <=( a3006a ) or ( a3001a );
 a3008a <=( a3007a ) or ( a2998a );
 a3011a <=( a1958a ) or ( a1959a );
 a3014a <=( a1956a ) or ( a1957a );
 a3015a <=( a3014a ) or ( a3011a );
 a3018a <=( a1954a ) or ( a1955a );
 a3022a <=( a1951a ) or ( a1952a );
 a3023a <=( a1953a ) or ( a3022a );
 a3024a <=( a3023a ) or ( a3018a );
 a3025a <=( a3024a ) or ( a3015a );
 a3026a <=( a3025a ) or ( a3008a );
 a3027a <=( a3026a ) or ( a2991a );
 a3028a <=( a3027a ) or ( a2956a );
 a3031a <=( a1949a ) or ( a1950a );
 a3034a <=( a1947a ) or ( a1948a );
 a3035a <=( a3034a ) or ( a3031a );
 a3038a <=( a1945a ) or ( a1946a );
 a3042a <=( a1942a ) or ( a1943a );
 a3043a <=( a1944a ) or ( a3042a );
 a3044a <=( a3043a ) or ( a3038a );
 a3045a <=( a3044a ) or ( a3035a );
 a3048a <=( a1940a ) or ( a1941a );
 a3051a <=( a1938a ) or ( a1939a );
 a3052a <=( a3051a ) or ( a3048a );
 a3055a <=( a1936a ) or ( a1937a );
 a3059a <=( a1933a ) or ( a1934a );
 a3060a <=( a1935a ) or ( a3059a );
 a3061a <=( a3060a ) or ( a3055a );
 a3062a <=( a3061a ) or ( a3052a );
 a3063a <=( a3062a ) or ( a3045a );
 a3066a <=( a1931a ) or ( a1932a );
 a3069a <=( a1929a ) or ( a1930a );
 a3070a <=( a3069a ) or ( a3066a );
 a3073a <=( a1927a ) or ( a1928a );
 a3077a <=( a1924a ) or ( a1925a );
 a3078a <=( a1926a ) or ( a3077a );
 a3079a <=( a3078a ) or ( a3073a );
 a3080a <=( a3079a ) or ( a3070a );
 a3083a <=( a1922a ) or ( a1923a );
 a3086a <=( a1920a ) or ( a1921a );
 a3087a <=( a3086a ) or ( a3083a );
 a3090a <=( a1918a ) or ( a1919a );
 a3094a <=( a1915a ) or ( a1916a );
 a3095a <=( a1917a ) or ( a3094a );
 a3096a <=( a3095a ) or ( a3090a );
 a3097a <=( a3096a ) or ( a3087a );
 a3098a <=( a3097a ) or ( a3080a );
 a3099a <=( a3098a ) or ( a3063a );
 a3102a <=( a1913a ) or ( a1914a );
 a3105a <=( a1911a ) or ( a1912a );
 a3106a <=( a3105a ) or ( a3102a );
 a3109a <=( a1909a ) or ( a1910a );
 a3113a <=( a1906a ) or ( a1907a );
 a3114a <=( a1908a ) or ( a3113a );
 a3115a <=( a3114a ) or ( a3109a );
 a3116a <=( a3115a ) or ( a3106a );
 a3119a <=( a1904a ) or ( a1905a );
 a3122a <=( a1902a ) or ( a1903a );
 a3123a <=( a3122a ) or ( a3119a );
 a3126a <=( a1900a ) or ( a1901a );
 a3130a <=( a1897a ) or ( a1898a );
 a3131a <=( a1899a ) or ( a3130a );
 a3132a <=( a3131a ) or ( a3126a );
 a3133a <=( a3132a ) or ( a3123a );
 a3134a <=( a3133a ) or ( a3116a );
 a3137a <=( a1895a ) or ( a1896a );
 a3140a <=( a1893a ) or ( a1894a );
 a3141a <=( a3140a ) or ( a3137a );
 a3144a <=( a1891a ) or ( a1892a );
 a3148a <=( a1888a ) or ( a1889a );
 a3149a <=( a1890a ) or ( a3148a );
 a3150a <=( a3149a ) or ( a3144a );
 a3151a <=( a3150a ) or ( a3141a );
 a3154a <=( a1886a ) or ( a1887a );
 a3157a <=( a1884a ) or ( a1885a );
 a3158a <=( a3157a ) or ( a3154a );
 a3161a <=( a1882a ) or ( a1883a );
 a3165a <=( a1879a ) or ( a1880a );
 a3166a <=( a1881a ) or ( a3165a );
 a3167a <=( a3166a ) or ( a3161a );
 a3168a <=( a3167a ) or ( a3158a );
 a3169a <=( a3168a ) or ( a3151a );
 a3170a <=( a3169a ) or ( a3134a );
 a3171a <=( a3170a ) or ( a3099a );
 a3172a <=( a3171a ) or ( a3028a );
 a3175a <=( a1877a ) or ( a1878a );
 a3178a <=( a1875a ) or ( a1876a );
 a3179a <=( a3178a ) or ( a3175a );
 a3182a <=( a1873a ) or ( a1874a );
 a3186a <=( a1870a ) or ( a1871a );
 a3187a <=( a1872a ) or ( a3186a );
 a3188a <=( a3187a ) or ( a3182a );
 a3189a <=( a3188a ) or ( a3179a );
 a3192a <=( a1868a ) or ( a1869a );
 a3195a <=( a1866a ) or ( a1867a );
 a3196a <=( a3195a ) or ( a3192a );
 a3199a <=( a1864a ) or ( a1865a );
 a3203a <=( a1861a ) or ( a1862a );
 a3204a <=( a1863a ) or ( a3203a );
 a3205a <=( a3204a ) or ( a3199a );
 a3206a <=( a3205a ) or ( a3196a );
 a3207a <=( a3206a ) or ( a3189a );
 a3210a <=( a1859a ) or ( a1860a );
 a3213a <=( a1857a ) or ( a1858a );
 a3214a <=( a3213a ) or ( a3210a );
 a3217a <=( a1855a ) or ( a1856a );
 a3221a <=( a1852a ) or ( a1853a );
 a3222a <=( a1854a ) or ( a3221a );
 a3223a <=( a3222a ) or ( a3217a );
 a3224a <=( a3223a ) or ( a3214a );
 a3227a <=( a1850a ) or ( a1851a );
 a3230a <=( a1848a ) or ( a1849a );
 a3231a <=( a3230a ) or ( a3227a );
 a3234a <=( a1846a ) or ( a1847a );
 a3238a <=( a1843a ) or ( a1844a );
 a3239a <=( a1845a ) or ( a3238a );
 a3240a <=( a3239a ) or ( a3234a );
 a3241a <=( a3240a ) or ( a3231a );
 a3242a <=( a3241a ) or ( a3224a );
 a3243a <=( a3242a ) or ( a3207a );
 a3246a <=( a1841a ) or ( a1842a );
 a3249a <=( a1839a ) or ( a1840a );
 a3250a <=( a3249a ) or ( a3246a );
 a3253a <=( a1837a ) or ( a1838a );
 a3257a <=( a1834a ) or ( a1835a );
 a3258a <=( a1836a ) or ( a3257a );
 a3259a <=( a3258a ) or ( a3253a );
 a3260a <=( a3259a ) or ( a3250a );
 a3263a <=( a1832a ) or ( a1833a );
 a3266a <=( a1830a ) or ( a1831a );
 a3267a <=( a3266a ) or ( a3263a );
 a3270a <=( a1828a ) or ( a1829a );
 a3274a <=( a1825a ) or ( a1826a );
 a3275a <=( a1827a ) or ( a3274a );
 a3276a <=( a3275a ) or ( a3270a );
 a3277a <=( a3276a ) or ( a3267a );
 a3278a <=( a3277a ) or ( a3260a );
 a3281a <=( a1823a ) or ( a1824a );
 a3284a <=( a1821a ) or ( a1822a );
 a3285a <=( a3284a ) or ( a3281a );
 a3288a <=( a1819a ) or ( a1820a );
 a3292a <=( a1816a ) or ( a1817a );
 a3293a <=( a1818a ) or ( a3292a );
 a3294a <=( a3293a ) or ( a3288a );
 a3295a <=( a3294a ) or ( a3285a );
 a3298a <=( a1814a ) or ( a1815a );
 a3301a <=( a1812a ) or ( a1813a );
 a3302a <=( a3301a ) or ( a3298a );
 a3305a <=( a1810a ) or ( a1811a );
 a3309a <=( a1807a ) or ( a1808a );
 a3310a <=( a1809a ) or ( a3309a );
 a3311a <=( a3310a ) or ( a3305a );
 a3312a <=( a3311a ) or ( a3302a );
 a3313a <=( a3312a ) or ( a3295a );
 a3314a <=( a3313a ) or ( a3278a );
 a3315a <=( a3314a ) or ( a3243a );
 a3318a <=( a1805a ) or ( a1806a );
 a3321a <=( a1803a ) or ( a1804a );
 a3322a <=( a3321a ) or ( a3318a );
 a3325a <=( a1801a ) or ( a1802a );
 a3329a <=( a1798a ) or ( a1799a );
 a3330a <=( a1800a ) or ( a3329a );
 a3331a <=( a3330a ) or ( a3325a );
 a3332a <=( a3331a ) or ( a3322a );
 a3335a <=( a1796a ) or ( a1797a );
 a3338a <=( a1794a ) or ( a1795a );
 a3339a <=( a3338a ) or ( a3335a );
 a3342a <=( a1792a ) or ( a1793a );
 a3346a <=( a1789a ) or ( a1790a );
 a3347a <=( a1791a ) or ( a3346a );
 a3348a <=( a3347a ) or ( a3342a );
 a3349a <=( a3348a ) or ( a3339a );
 a3350a <=( a3349a ) or ( a3332a );
 a3353a <=( a1787a ) or ( a1788a );
 a3356a <=( a1785a ) or ( a1786a );
 a3357a <=( a3356a ) or ( a3353a );
 a3360a <=( a1783a ) or ( a1784a );
 a3364a <=( a1780a ) or ( a1781a );
 a3365a <=( a1782a ) or ( a3364a );
 a3366a <=( a3365a ) or ( a3360a );
 a3367a <=( a3366a ) or ( a3357a );
 a3370a <=( a1778a ) or ( a1779a );
 a3373a <=( a1776a ) or ( a1777a );
 a3374a <=( a3373a ) or ( a3370a );
 a3377a <=( a1774a ) or ( a1775a );
 a3381a <=( a1771a ) or ( a1772a );
 a3382a <=( a1773a ) or ( a3381a );
 a3383a <=( a3382a ) or ( a3377a );
 a3384a <=( a3383a ) or ( a3374a );
 a3385a <=( a3384a ) or ( a3367a );
 a3386a <=( a3385a ) or ( a3350a );
 a3389a <=( a1769a ) or ( a1770a );
 a3392a <=( a1767a ) or ( a1768a );
 a3393a <=( a3392a ) or ( a3389a );
 a3396a <=( a1765a ) or ( a1766a );
 a3400a <=( a1762a ) or ( a1763a );
 a3401a <=( a1764a ) or ( a3400a );
 a3402a <=( a3401a ) or ( a3396a );
 a3403a <=( a3402a ) or ( a3393a );
 a3406a <=( a1760a ) or ( a1761a );
 a3409a <=( a1758a ) or ( a1759a );
 a3410a <=( a3409a ) or ( a3406a );
 a3413a <=( a1756a ) or ( a1757a );
 a3417a <=( a1753a ) or ( a1754a );
 a3418a <=( a1755a ) or ( a3417a );
 a3419a <=( a3418a ) or ( a3413a );
 a3420a <=( a3419a ) or ( a3410a );
 a3421a <=( a3420a ) or ( a3403a );
 a3424a <=( a1751a ) or ( a1752a );
 a3427a <=( a1749a ) or ( a1750a );
 a3428a <=( a3427a ) or ( a3424a );
 a3431a <=( a1747a ) or ( a1748a );
 a3435a <=( a1744a ) or ( a1745a );
 a3436a <=( a1746a ) or ( a3435a );
 a3437a <=( a3436a ) or ( a3431a );
 a3438a <=( a3437a ) or ( a3428a );
 a3441a <=( a1742a ) or ( a1743a );
 a3445a <=( a1739a ) or ( a1740a );
 a3446a <=( a1741a ) or ( a3445a );
 a3447a <=( a3446a ) or ( a3441a );
 a3450a <=( a1737a ) or ( a1738a );
 a3454a <=( a1734a ) or ( a1735a );
 a3455a <=( a1736a ) or ( a3454a );
 a3456a <=( a3455a ) or ( a3450a );
 a3457a <=( a3456a ) or ( a3447a );
 a3458a <=( a3457a ) or ( a3438a );
 a3459a <=( a3458a ) or ( a3421a );
 a3460a <=( a3459a ) or ( a3386a );
 a3461a <=( a3460a ) or ( a3315a );
 a3462a <=( a3461a ) or ( a3172a );
 a3463a <=( a3462a ) or ( a2885a );
 a3466a <=( a1732a ) or ( a1733a );
 a3469a <=( a1730a ) or ( a1731a );
 a3470a <=( a3469a ) or ( a3466a );
 a3473a <=( a1728a ) or ( a1729a );
 a3477a <=( a1725a ) or ( a1726a );
 a3478a <=( a1727a ) or ( a3477a );
 a3479a <=( a3478a ) or ( a3473a );
 a3480a <=( a3479a ) or ( a3470a );
 a3483a <=( a1723a ) or ( a1724a );
 a3486a <=( a1721a ) or ( a1722a );
 a3487a <=( a3486a ) or ( a3483a );
 a3490a <=( a1719a ) or ( a1720a );
 a3494a <=( a1716a ) or ( a1717a );
 a3495a <=( a1718a ) or ( a3494a );
 a3496a <=( a3495a ) or ( a3490a );
 a3497a <=( a3496a ) or ( a3487a );
 a3498a <=( a3497a ) or ( a3480a );
 a3501a <=( a1714a ) or ( a1715a );
 a3504a <=( a1712a ) or ( a1713a );
 a3505a <=( a3504a ) or ( a3501a );
 a3508a <=( a1710a ) or ( a1711a );
 a3512a <=( a1707a ) or ( a1708a );
 a3513a <=( a1709a ) or ( a3512a );
 a3514a <=( a3513a ) or ( a3508a );
 a3515a <=( a3514a ) or ( a3505a );
 a3518a <=( a1705a ) or ( a1706a );
 a3521a <=( a1703a ) or ( a1704a );
 a3522a <=( a3521a ) or ( a3518a );
 a3525a <=( a1701a ) or ( a1702a );
 a3529a <=( a1698a ) or ( a1699a );
 a3530a <=( a1700a ) or ( a3529a );
 a3531a <=( a3530a ) or ( a3525a );
 a3532a <=( a3531a ) or ( a3522a );
 a3533a <=( a3532a ) or ( a3515a );
 a3534a <=( a3533a ) or ( a3498a );
 a3537a <=( a1696a ) or ( a1697a );
 a3540a <=( a1694a ) or ( a1695a );
 a3541a <=( a3540a ) or ( a3537a );
 a3544a <=( a1692a ) or ( a1693a );
 a3548a <=( a1689a ) or ( a1690a );
 a3549a <=( a1691a ) or ( a3548a );
 a3550a <=( a3549a ) or ( a3544a );
 a3551a <=( a3550a ) or ( a3541a );
 a3554a <=( a1687a ) or ( a1688a );
 a3557a <=( a1685a ) or ( a1686a );
 a3558a <=( a3557a ) or ( a3554a );
 a3561a <=( a1683a ) or ( a1684a );
 a3565a <=( a1680a ) or ( a1681a );
 a3566a <=( a1682a ) or ( a3565a );
 a3567a <=( a3566a ) or ( a3561a );
 a3568a <=( a3567a ) or ( a3558a );
 a3569a <=( a3568a ) or ( a3551a );
 a3572a <=( a1678a ) or ( a1679a );
 a3575a <=( a1676a ) or ( a1677a );
 a3576a <=( a3575a ) or ( a3572a );
 a3579a <=( a1674a ) or ( a1675a );
 a3583a <=( a1671a ) or ( a1672a );
 a3584a <=( a1673a ) or ( a3583a );
 a3585a <=( a3584a ) or ( a3579a );
 a3586a <=( a3585a ) or ( a3576a );
 a3589a <=( a1669a ) or ( a1670a );
 a3592a <=( a1667a ) or ( a1668a );
 a3593a <=( a3592a ) or ( a3589a );
 a3596a <=( a1665a ) or ( a1666a );
 a3600a <=( a1662a ) or ( a1663a );
 a3601a <=( a1664a ) or ( a3600a );
 a3602a <=( a3601a ) or ( a3596a );
 a3603a <=( a3602a ) or ( a3593a );
 a3604a <=( a3603a ) or ( a3586a );
 a3605a <=( a3604a ) or ( a3569a );
 a3606a <=( a3605a ) or ( a3534a );
 a3609a <=( a1660a ) or ( a1661a );
 a3612a <=( a1658a ) or ( a1659a );
 a3613a <=( a3612a ) or ( a3609a );
 a3616a <=( a1656a ) or ( a1657a );
 a3620a <=( a1653a ) or ( a1654a );
 a3621a <=( a1655a ) or ( a3620a );
 a3622a <=( a3621a ) or ( a3616a );
 a3623a <=( a3622a ) or ( a3613a );
 a3626a <=( a1651a ) or ( a1652a );
 a3629a <=( a1649a ) or ( a1650a );
 a3630a <=( a3629a ) or ( a3626a );
 a3633a <=( a1647a ) or ( a1648a );
 a3637a <=( a1644a ) or ( a1645a );
 a3638a <=( a1646a ) or ( a3637a );
 a3639a <=( a3638a ) or ( a3633a );
 a3640a <=( a3639a ) or ( a3630a );
 a3641a <=( a3640a ) or ( a3623a );
 a3644a <=( a1642a ) or ( a1643a );
 a3647a <=( a1640a ) or ( a1641a );
 a3648a <=( a3647a ) or ( a3644a );
 a3651a <=( a1638a ) or ( a1639a );
 a3655a <=( a1635a ) or ( a1636a );
 a3656a <=( a1637a ) or ( a3655a );
 a3657a <=( a3656a ) or ( a3651a );
 a3658a <=( a3657a ) or ( a3648a );
 a3661a <=( a1633a ) or ( a1634a );
 a3664a <=( a1631a ) or ( a1632a );
 a3665a <=( a3664a ) or ( a3661a );
 a3668a <=( a1629a ) or ( a1630a );
 a3672a <=( a1626a ) or ( a1627a );
 a3673a <=( a1628a ) or ( a3672a );
 a3674a <=( a3673a ) or ( a3668a );
 a3675a <=( a3674a ) or ( a3665a );
 a3676a <=( a3675a ) or ( a3658a );
 a3677a <=( a3676a ) or ( a3641a );
 a3680a <=( a1624a ) or ( a1625a );
 a3683a <=( a1622a ) or ( a1623a );
 a3684a <=( a3683a ) or ( a3680a );
 a3687a <=( a1620a ) or ( a1621a );
 a3691a <=( a1617a ) or ( a1618a );
 a3692a <=( a1619a ) or ( a3691a );
 a3693a <=( a3692a ) or ( a3687a );
 a3694a <=( a3693a ) or ( a3684a );
 a3697a <=( a1615a ) or ( a1616a );
 a3700a <=( a1613a ) or ( a1614a );
 a3701a <=( a3700a ) or ( a3697a );
 a3704a <=( a1611a ) or ( a1612a );
 a3708a <=( a1608a ) or ( a1609a );
 a3709a <=( a1610a ) or ( a3708a );
 a3710a <=( a3709a ) or ( a3704a );
 a3711a <=( a3710a ) or ( a3701a );
 a3712a <=( a3711a ) or ( a3694a );
 a3715a <=( a1606a ) or ( a1607a );
 a3718a <=( a1604a ) or ( a1605a );
 a3719a <=( a3718a ) or ( a3715a );
 a3722a <=( a1602a ) or ( a1603a );
 a3726a <=( a1599a ) or ( a1600a );
 a3727a <=( a1601a ) or ( a3726a );
 a3728a <=( a3727a ) or ( a3722a );
 a3729a <=( a3728a ) or ( a3719a );
 a3732a <=( a1597a ) or ( a1598a );
 a3735a <=( a1595a ) or ( a1596a );
 a3736a <=( a3735a ) or ( a3732a );
 a3739a <=( a1593a ) or ( a1594a );
 a3743a <=( a1590a ) or ( a1591a );
 a3744a <=( a1592a ) or ( a3743a );
 a3745a <=( a3744a ) or ( a3739a );
 a3746a <=( a3745a ) or ( a3736a );
 a3747a <=( a3746a ) or ( a3729a );
 a3748a <=( a3747a ) or ( a3712a );
 a3749a <=( a3748a ) or ( a3677a );
 a3750a <=( a3749a ) or ( a3606a );
 a3753a <=( a1588a ) or ( a1589a );
 a3756a <=( a1586a ) or ( a1587a );
 a3757a <=( a3756a ) or ( a3753a );
 a3760a <=( a1584a ) or ( a1585a );
 a3764a <=( a1581a ) or ( a1582a );
 a3765a <=( a1583a ) or ( a3764a );
 a3766a <=( a3765a ) or ( a3760a );
 a3767a <=( a3766a ) or ( a3757a );
 a3770a <=( a1579a ) or ( a1580a );
 a3773a <=( a1577a ) or ( a1578a );
 a3774a <=( a3773a ) or ( a3770a );
 a3777a <=( a1575a ) or ( a1576a );
 a3781a <=( a1572a ) or ( a1573a );
 a3782a <=( a1574a ) or ( a3781a );
 a3783a <=( a3782a ) or ( a3777a );
 a3784a <=( a3783a ) or ( a3774a );
 a3785a <=( a3784a ) or ( a3767a );
 a3788a <=( a1570a ) or ( a1571a );
 a3791a <=( a1568a ) or ( a1569a );
 a3792a <=( a3791a ) or ( a3788a );
 a3795a <=( a1566a ) or ( a1567a );
 a3799a <=( a1563a ) or ( a1564a );
 a3800a <=( a1565a ) or ( a3799a );
 a3801a <=( a3800a ) or ( a3795a );
 a3802a <=( a3801a ) or ( a3792a );
 a3805a <=( a1561a ) or ( a1562a );
 a3808a <=( a1559a ) or ( a1560a );
 a3809a <=( a3808a ) or ( a3805a );
 a3812a <=( a1557a ) or ( a1558a );
 a3816a <=( a1554a ) or ( a1555a );
 a3817a <=( a1556a ) or ( a3816a );
 a3818a <=( a3817a ) or ( a3812a );
 a3819a <=( a3818a ) or ( a3809a );
 a3820a <=( a3819a ) or ( a3802a );
 a3821a <=( a3820a ) or ( a3785a );
 a3824a <=( a1552a ) or ( a1553a );
 a3827a <=( a1550a ) or ( a1551a );
 a3828a <=( a3827a ) or ( a3824a );
 a3831a <=( a1548a ) or ( a1549a );
 a3835a <=( a1545a ) or ( a1546a );
 a3836a <=( a1547a ) or ( a3835a );
 a3837a <=( a3836a ) or ( a3831a );
 a3838a <=( a3837a ) or ( a3828a );
 a3841a <=( a1543a ) or ( a1544a );
 a3844a <=( a1541a ) or ( a1542a );
 a3845a <=( a3844a ) or ( a3841a );
 a3848a <=( a1539a ) or ( a1540a );
 a3852a <=( a1536a ) or ( a1537a );
 a3853a <=( a1538a ) or ( a3852a );
 a3854a <=( a3853a ) or ( a3848a );
 a3855a <=( a3854a ) or ( a3845a );
 a3856a <=( a3855a ) or ( a3838a );
 a3859a <=( a1534a ) or ( a1535a );
 a3862a <=( a1532a ) or ( a1533a );
 a3863a <=( a3862a ) or ( a3859a );
 a3866a <=( a1530a ) or ( a1531a );
 a3870a <=( a1527a ) or ( a1528a );
 a3871a <=( a1529a ) or ( a3870a );
 a3872a <=( a3871a ) or ( a3866a );
 a3873a <=( a3872a ) or ( a3863a );
 a3876a <=( a1525a ) or ( a1526a );
 a3879a <=( a1523a ) or ( a1524a );
 a3880a <=( a3879a ) or ( a3876a );
 a3883a <=( a1521a ) or ( a1522a );
 a3887a <=( a1518a ) or ( a1519a );
 a3888a <=( a1520a ) or ( a3887a );
 a3889a <=( a3888a ) or ( a3883a );
 a3890a <=( a3889a ) or ( a3880a );
 a3891a <=( a3890a ) or ( a3873a );
 a3892a <=( a3891a ) or ( a3856a );
 a3893a <=( a3892a ) or ( a3821a );
 a3896a <=( a1516a ) or ( a1517a );
 a3899a <=( a1514a ) or ( a1515a );
 a3900a <=( a3899a ) or ( a3896a );
 a3903a <=( a1512a ) or ( a1513a );
 a3907a <=( a1509a ) or ( a1510a );
 a3908a <=( a1511a ) or ( a3907a );
 a3909a <=( a3908a ) or ( a3903a );
 a3910a <=( a3909a ) or ( a3900a );
 a3913a <=( a1507a ) or ( a1508a );
 a3916a <=( a1505a ) or ( a1506a );
 a3917a <=( a3916a ) or ( a3913a );
 a3920a <=( a1503a ) or ( a1504a );
 a3924a <=( a1500a ) or ( a1501a );
 a3925a <=( a1502a ) or ( a3924a );
 a3926a <=( a3925a ) or ( a3920a );
 a3927a <=( a3926a ) or ( a3917a );
 a3928a <=( a3927a ) or ( a3910a );
 a3931a <=( a1498a ) or ( a1499a );
 a3934a <=( a1496a ) or ( a1497a );
 a3935a <=( a3934a ) or ( a3931a );
 a3938a <=( a1494a ) or ( a1495a );
 a3942a <=( a1491a ) or ( a1492a );
 a3943a <=( a1493a ) or ( a3942a );
 a3944a <=( a3943a ) or ( a3938a );
 a3945a <=( a3944a ) or ( a3935a );
 a3948a <=( a1489a ) or ( a1490a );
 a3951a <=( a1487a ) or ( a1488a );
 a3952a <=( a3951a ) or ( a3948a );
 a3955a <=( a1485a ) or ( a1486a );
 a3959a <=( a1482a ) or ( a1483a );
 a3960a <=( a1484a ) or ( a3959a );
 a3961a <=( a3960a ) or ( a3955a );
 a3962a <=( a3961a ) or ( a3952a );
 a3963a <=( a3962a ) or ( a3945a );
 a3964a <=( a3963a ) or ( a3928a );
 a3967a <=( a1480a ) or ( a1481a );
 a3970a <=( a1478a ) or ( a1479a );
 a3971a <=( a3970a ) or ( a3967a );
 a3974a <=( a1476a ) or ( a1477a );
 a3978a <=( a1473a ) or ( a1474a );
 a3979a <=( a1475a ) or ( a3978a );
 a3980a <=( a3979a ) or ( a3974a );
 a3981a <=( a3980a ) or ( a3971a );
 a3984a <=( a1471a ) or ( a1472a );
 a3987a <=( a1469a ) or ( a1470a );
 a3988a <=( a3987a ) or ( a3984a );
 a3991a <=( a1467a ) or ( a1468a );
 a3995a <=( a1464a ) or ( a1465a );
 a3996a <=( a1466a ) or ( a3995a );
 a3997a <=( a3996a ) or ( a3991a );
 a3998a <=( a3997a ) or ( a3988a );
 a3999a <=( a3998a ) or ( a3981a );
 a4002a <=( a1462a ) or ( a1463a );
 a4005a <=( a1460a ) or ( a1461a );
 a4006a <=( a4005a ) or ( a4002a );
 a4009a <=( a1458a ) or ( a1459a );
 a4013a <=( a1455a ) or ( a1456a );
 a4014a <=( a1457a ) or ( a4013a );
 a4015a <=( a4014a ) or ( a4009a );
 a4016a <=( a4015a ) or ( a4006a );
 a4019a <=( a1453a ) or ( a1454a );
 a4023a <=( a1450a ) or ( a1451a );
 a4024a <=( a1452a ) or ( a4023a );
 a4025a <=( a4024a ) or ( a4019a );
 a4028a <=( a1448a ) or ( a1449a );
 a4032a <=( a1445a ) or ( a1446a );
 a4033a <=( a1447a ) or ( a4032a );
 a4034a <=( a4033a ) or ( a4028a );
 a4035a <=( a4034a ) or ( a4025a );
 a4036a <=( a4035a ) or ( a4016a );
 a4037a <=( a4036a ) or ( a3999a );
 a4038a <=( a4037a ) or ( a3964a );
 a4039a <=( a4038a ) or ( a3893a );
 a4040a <=( a4039a ) or ( a3750a );
 a4043a <=( a1443a ) or ( a1444a );
 a4046a <=( a1441a ) or ( a1442a );
 a4047a <=( a4046a ) or ( a4043a );
 a4050a <=( a1439a ) or ( a1440a );
 a4054a <=( a1436a ) or ( a1437a );
 a4055a <=( a1438a ) or ( a4054a );
 a4056a <=( a4055a ) or ( a4050a );
 a4057a <=( a4056a ) or ( a4047a );
 a4060a <=( a1434a ) or ( a1435a );
 a4063a <=( a1432a ) or ( a1433a );
 a4064a <=( a4063a ) or ( a4060a );
 a4067a <=( a1430a ) or ( a1431a );
 a4071a <=( a1427a ) or ( a1428a );
 a4072a <=( a1429a ) or ( a4071a );
 a4073a <=( a4072a ) or ( a4067a );
 a4074a <=( a4073a ) or ( a4064a );
 a4075a <=( a4074a ) or ( a4057a );
 a4078a <=( a1425a ) or ( a1426a );
 a4081a <=( a1423a ) or ( a1424a );
 a4082a <=( a4081a ) or ( a4078a );
 a4085a <=( a1421a ) or ( a1422a );
 a4089a <=( a1418a ) or ( a1419a );
 a4090a <=( a1420a ) or ( a4089a );
 a4091a <=( a4090a ) or ( a4085a );
 a4092a <=( a4091a ) or ( a4082a );
 a4095a <=( a1416a ) or ( a1417a );
 a4098a <=( a1414a ) or ( a1415a );
 a4099a <=( a4098a ) or ( a4095a );
 a4102a <=( a1412a ) or ( a1413a );
 a4106a <=( a1409a ) or ( a1410a );
 a4107a <=( a1411a ) or ( a4106a );
 a4108a <=( a4107a ) or ( a4102a );
 a4109a <=( a4108a ) or ( a4099a );
 a4110a <=( a4109a ) or ( a4092a );
 a4111a <=( a4110a ) or ( a4075a );
 a4114a <=( a1407a ) or ( a1408a );
 a4117a <=( a1405a ) or ( a1406a );
 a4118a <=( a4117a ) or ( a4114a );
 a4121a <=( a1403a ) or ( a1404a );
 a4125a <=( a1400a ) or ( a1401a );
 a4126a <=( a1402a ) or ( a4125a );
 a4127a <=( a4126a ) or ( a4121a );
 a4128a <=( a4127a ) or ( a4118a );
 a4131a <=( a1398a ) or ( a1399a );
 a4134a <=( a1396a ) or ( a1397a );
 a4135a <=( a4134a ) or ( a4131a );
 a4138a <=( a1394a ) or ( a1395a );
 a4142a <=( a1391a ) or ( a1392a );
 a4143a <=( a1393a ) or ( a4142a );
 a4144a <=( a4143a ) or ( a4138a );
 a4145a <=( a4144a ) or ( a4135a );
 a4146a <=( a4145a ) or ( a4128a );
 a4149a <=( a1389a ) or ( a1390a );
 a4152a <=( a1387a ) or ( a1388a );
 a4153a <=( a4152a ) or ( a4149a );
 a4156a <=( a1385a ) or ( a1386a );
 a4160a <=( a1382a ) or ( a1383a );
 a4161a <=( a1384a ) or ( a4160a );
 a4162a <=( a4161a ) or ( a4156a );
 a4163a <=( a4162a ) or ( a4153a );
 a4166a <=( a1380a ) or ( a1381a );
 a4169a <=( a1378a ) or ( a1379a );
 a4170a <=( a4169a ) or ( a4166a );
 a4173a <=( a1376a ) or ( a1377a );
 a4177a <=( a1373a ) or ( a1374a );
 a4178a <=( a1375a ) or ( a4177a );
 a4179a <=( a4178a ) or ( a4173a );
 a4180a <=( a4179a ) or ( a4170a );
 a4181a <=( a4180a ) or ( a4163a );
 a4182a <=( a4181a ) or ( a4146a );
 a4183a <=( a4182a ) or ( a4111a );
 a4186a <=( a1371a ) or ( a1372a );
 a4189a <=( a1369a ) or ( a1370a );
 a4190a <=( a4189a ) or ( a4186a );
 a4193a <=( a1367a ) or ( a1368a );
 a4197a <=( a1364a ) or ( a1365a );
 a4198a <=( a1366a ) or ( a4197a );
 a4199a <=( a4198a ) or ( a4193a );
 a4200a <=( a4199a ) or ( a4190a );
 a4203a <=( a1362a ) or ( a1363a );
 a4206a <=( a1360a ) or ( a1361a );
 a4207a <=( a4206a ) or ( a4203a );
 a4210a <=( a1358a ) or ( a1359a );
 a4214a <=( a1355a ) or ( a1356a );
 a4215a <=( a1357a ) or ( a4214a );
 a4216a <=( a4215a ) or ( a4210a );
 a4217a <=( a4216a ) or ( a4207a );
 a4218a <=( a4217a ) or ( a4200a );
 a4221a <=( a1353a ) or ( a1354a );
 a4224a <=( a1351a ) or ( a1352a );
 a4225a <=( a4224a ) or ( a4221a );
 a4228a <=( a1349a ) or ( a1350a );
 a4232a <=( a1346a ) or ( a1347a );
 a4233a <=( a1348a ) or ( a4232a );
 a4234a <=( a4233a ) or ( a4228a );
 a4235a <=( a4234a ) or ( a4225a );
 a4238a <=( a1344a ) or ( a1345a );
 a4241a <=( a1342a ) or ( a1343a );
 a4242a <=( a4241a ) or ( a4238a );
 a4245a <=( a1340a ) or ( a1341a );
 a4249a <=( a1337a ) or ( a1338a );
 a4250a <=( a1339a ) or ( a4249a );
 a4251a <=( a4250a ) or ( a4245a );
 a4252a <=( a4251a ) or ( a4242a );
 a4253a <=( a4252a ) or ( a4235a );
 a4254a <=( a4253a ) or ( a4218a );
 a4257a <=( a1335a ) or ( a1336a );
 a4260a <=( a1333a ) or ( a1334a );
 a4261a <=( a4260a ) or ( a4257a );
 a4264a <=( a1331a ) or ( a1332a );
 a4268a <=( a1328a ) or ( a1329a );
 a4269a <=( a1330a ) or ( a4268a );
 a4270a <=( a4269a ) or ( a4264a );
 a4271a <=( a4270a ) or ( a4261a );
 a4274a <=( a1326a ) or ( a1327a );
 a4277a <=( a1324a ) or ( a1325a );
 a4278a <=( a4277a ) or ( a4274a );
 a4281a <=( a1322a ) or ( a1323a );
 a4285a <=( a1319a ) or ( a1320a );
 a4286a <=( a1321a ) or ( a4285a );
 a4287a <=( a4286a ) or ( a4281a );
 a4288a <=( a4287a ) or ( a4278a );
 a4289a <=( a4288a ) or ( a4271a );
 a4292a <=( a1317a ) or ( a1318a );
 a4295a <=( a1315a ) or ( a1316a );
 a4296a <=( a4295a ) or ( a4292a );
 a4299a <=( a1313a ) or ( a1314a );
 a4303a <=( a1310a ) or ( a1311a );
 a4304a <=( a1312a ) or ( a4303a );
 a4305a <=( a4304a ) or ( a4299a );
 a4306a <=( a4305a ) or ( a4296a );
 a4309a <=( a1308a ) or ( a1309a );
 a4312a <=( a1306a ) or ( a1307a );
 a4313a <=( a4312a ) or ( a4309a );
 a4316a <=( a1304a ) or ( a1305a );
 a4320a <=( a1301a ) or ( a1302a );
 a4321a <=( a1303a ) or ( a4320a );
 a4322a <=( a4321a ) or ( a4316a );
 a4323a <=( a4322a ) or ( a4313a );
 a4324a <=( a4323a ) or ( a4306a );
 a4325a <=( a4324a ) or ( a4289a );
 a4326a <=( a4325a ) or ( a4254a );
 a4327a <=( a4326a ) or ( a4183a );
 a4330a <=( a1299a ) or ( a1300a );
 a4333a <=( a1297a ) or ( a1298a );
 a4334a <=( a4333a ) or ( a4330a );
 a4337a <=( a1295a ) or ( a1296a );
 a4341a <=( a1292a ) or ( a1293a );
 a4342a <=( a1294a ) or ( a4341a );
 a4343a <=( a4342a ) or ( a4337a );
 a4344a <=( a4343a ) or ( a4334a );
 a4347a <=( a1290a ) or ( a1291a );
 a4350a <=( a1288a ) or ( a1289a );
 a4351a <=( a4350a ) or ( a4347a );
 a4354a <=( a1286a ) or ( a1287a );
 a4358a <=( a1283a ) or ( a1284a );
 a4359a <=( a1285a ) or ( a4358a );
 a4360a <=( a4359a ) or ( a4354a );
 a4361a <=( a4360a ) or ( a4351a );
 a4362a <=( a4361a ) or ( a4344a );
 a4365a <=( a1281a ) or ( a1282a );
 a4368a <=( a1279a ) or ( a1280a );
 a4369a <=( a4368a ) or ( a4365a );
 a4372a <=( a1277a ) or ( a1278a );
 a4376a <=( a1274a ) or ( a1275a );
 a4377a <=( a1276a ) or ( a4376a );
 a4378a <=( a4377a ) or ( a4372a );
 a4379a <=( a4378a ) or ( a4369a );
 a4382a <=( a1272a ) or ( a1273a );
 a4385a <=( a1270a ) or ( a1271a );
 a4386a <=( a4385a ) or ( a4382a );
 a4389a <=( a1268a ) or ( a1269a );
 a4393a <=( a1265a ) or ( a1266a );
 a4394a <=( a1267a ) or ( a4393a );
 a4395a <=( a4394a ) or ( a4389a );
 a4396a <=( a4395a ) or ( a4386a );
 a4397a <=( a4396a ) or ( a4379a );
 a4398a <=( a4397a ) or ( a4362a );
 a4401a <=( a1263a ) or ( a1264a );
 a4404a <=( a1261a ) or ( a1262a );
 a4405a <=( a4404a ) or ( a4401a );
 a4408a <=( a1259a ) or ( a1260a );
 a4412a <=( a1256a ) or ( a1257a );
 a4413a <=( a1258a ) or ( a4412a );
 a4414a <=( a4413a ) or ( a4408a );
 a4415a <=( a4414a ) or ( a4405a );
 a4418a <=( a1254a ) or ( a1255a );
 a4421a <=( a1252a ) or ( a1253a );
 a4422a <=( a4421a ) or ( a4418a );
 a4425a <=( a1250a ) or ( a1251a );
 a4429a <=( a1247a ) or ( a1248a );
 a4430a <=( a1249a ) or ( a4429a );
 a4431a <=( a4430a ) or ( a4425a );
 a4432a <=( a4431a ) or ( a4422a );
 a4433a <=( a4432a ) or ( a4415a );
 a4436a <=( a1245a ) or ( a1246a );
 a4439a <=( a1243a ) or ( a1244a );
 a4440a <=( a4439a ) or ( a4436a );
 a4443a <=( a1241a ) or ( a1242a );
 a4447a <=( a1238a ) or ( a1239a );
 a4448a <=( a1240a ) or ( a4447a );
 a4449a <=( a4448a ) or ( a4443a );
 a4450a <=( a4449a ) or ( a4440a );
 a4453a <=( a1236a ) or ( a1237a );
 a4456a <=( a1234a ) or ( a1235a );
 a4457a <=( a4456a ) or ( a4453a );
 a4460a <=( a1232a ) or ( a1233a );
 a4464a <=( a1229a ) or ( a1230a );
 a4465a <=( a1231a ) or ( a4464a );
 a4466a <=( a4465a ) or ( a4460a );
 a4467a <=( a4466a ) or ( a4457a );
 a4468a <=( a4467a ) or ( a4450a );
 a4469a <=( a4468a ) or ( a4433a );
 a4470a <=( a4469a ) or ( a4398a );
 a4473a <=( a1227a ) or ( a1228a );
 a4476a <=( a1225a ) or ( a1226a );
 a4477a <=( a4476a ) or ( a4473a );
 a4480a <=( a1223a ) or ( a1224a );
 a4484a <=( a1220a ) or ( a1221a );
 a4485a <=( a1222a ) or ( a4484a );
 a4486a <=( a4485a ) or ( a4480a );
 a4487a <=( a4486a ) or ( a4477a );
 a4490a <=( a1218a ) or ( a1219a );
 a4493a <=( a1216a ) or ( a1217a );
 a4494a <=( a4493a ) or ( a4490a );
 a4497a <=( a1214a ) or ( a1215a );
 a4501a <=( a1211a ) or ( a1212a );
 a4502a <=( a1213a ) or ( a4501a );
 a4503a <=( a4502a ) or ( a4497a );
 a4504a <=( a4503a ) or ( a4494a );
 a4505a <=( a4504a ) or ( a4487a );
 a4508a <=( a1209a ) or ( a1210a );
 a4511a <=( a1207a ) or ( a1208a );
 a4512a <=( a4511a ) or ( a4508a );
 a4515a <=( a1205a ) or ( a1206a );
 a4519a <=( a1202a ) or ( a1203a );
 a4520a <=( a1204a ) or ( a4519a );
 a4521a <=( a4520a ) or ( a4515a );
 a4522a <=( a4521a ) or ( a4512a );
 a4525a <=( a1200a ) or ( a1201a );
 a4528a <=( a1198a ) or ( a1199a );
 a4529a <=( a4528a ) or ( a4525a );
 a4532a <=( a1196a ) or ( a1197a );
 a4536a <=( a1193a ) or ( a1194a );
 a4537a <=( a1195a ) or ( a4536a );
 a4538a <=( a4537a ) or ( a4532a );
 a4539a <=( a4538a ) or ( a4529a );
 a4540a <=( a4539a ) or ( a4522a );
 a4541a <=( a4540a ) or ( a4505a );
 a4544a <=( a1191a ) or ( a1192a );
 a4547a <=( a1189a ) or ( a1190a );
 a4548a <=( a4547a ) or ( a4544a );
 a4551a <=( a1187a ) or ( a1188a );
 a4555a <=( a1184a ) or ( a1185a );
 a4556a <=( a1186a ) or ( a4555a );
 a4557a <=( a4556a ) or ( a4551a );
 a4558a <=( a4557a ) or ( a4548a );
 a4561a <=( a1182a ) or ( a1183a );
 a4564a <=( a1180a ) or ( a1181a );
 a4565a <=( a4564a ) or ( a4561a );
 a4568a <=( a1178a ) or ( a1179a );
 a4572a <=( a1175a ) or ( a1176a );
 a4573a <=( a1177a ) or ( a4572a );
 a4574a <=( a4573a ) or ( a4568a );
 a4575a <=( a4574a ) or ( a4565a );
 a4576a <=( a4575a ) or ( a4558a );
 a4579a <=( a1173a ) or ( a1174a );
 a4582a <=( a1171a ) or ( a1172a );
 a4583a <=( a4582a ) or ( a4579a );
 a4586a <=( a1169a ) or ( a1170a );
 a4590a <=( a1166a ) or ( a1167a );
 a4591a <=( a1168a ) or ( a4590a );
 a4592a <=( a4591a ) or ( a4586a );
 a4593a <=( a4592a ) or ( a4583a );
 a4596a <=( a1164a ) or ( a1165a );
 a4600a <=( a1161a ) or ( a1162a );
 a4601a <=( a1163a ) or ( a4600a );
 a4602a <=( a4601a ) or ( a4596a );
 a4605a <=( a1159a ) or ( a1160a );
 a4609a <=( a1156a ) or ( a1157a );
 a4610a <=( a1158a ) or ( a4609a );
 a4611a <=( a4610a ) or ( a4605a );
 a4612a <=( a4611a ) or ( a4602a );
 a4613a <=( a4612a ) or ( a4593a );
 a4614a <=( a4613a ) or ( a4576a );
 a4615a <=( a4614a ) or ( a4541a );
 a4616a <=( a4615a ) or ( a4470a );
 a4617a <=( a4616a ) or ( a4327a );
 a4618a <=( a4617a ) or ( a4040a );
 a4619a <=( a4618a ) or ( a3463a );
 a4622a <=( a1154a ) or ( a1155a );
 a4625a <=( a1152a ) or ( a1153a );
 a4626a <=( a4625a ) or ( a4622a );
 a4629a <=( a1150a ) or ( a1151a );
 a4633a <=( a1147a ) or ( a1148a );
 a4634a <=( a1149a ) or ( a4633a );
 a4635a <=( a4634a ) or ( a4629a );
 a4636a <=( a4635a ) or ( a4626a );
 a4639a <=( a1145a ) or ( a1146a );
 a4642a <=( a1143a ) or ( a1144a );
 a4643a <=( a4642a ) or ( a4639a );
 a4646a <=( a1141a ) or ( a1142a );
 a4650a <=( a1138a ) or ( a1139a );
 a4651a <=( a1140a ) or ( a4650a );
 a4652a <=( a4651a ) or ( a4646a );
 a4653a <=( a4652a ) or ( a4643a );
 a4654a <=( a4653a ) or ( a4636a );
 a4657a <=( a1136a ) or ( a1137a );
 a4660a <=( a1134a ) or ( a1135a );
 a4661a <=( a4660a ) or ( a4657a );
 a4664a <=( a1132a ) or ( a1133a );
 a4668a <=( a1129a ) or ( a1130a );
 a4669a <=( a1131a ) or ( a4668a );
 a4670a <=( a4669a ) or ( a4664a );
 a4671a <=( a4670a ) or ( a4661a );
 a4674a <=( a1127a ) or ( a1128a );
 a4677a <=( a1125a ) or ( a1126a );
 a4678a <=( a4677a ) or ( a4674a );
 a4681a <=( a1123a ) or ( a1124a );
 a4685a <=( a1120a ) or ( a1121a );
 a4686a <=( a1122a ) or ( a4685a );
 a4687a <=( a4686a ) or ( a4681a );
 a4688a <=( a4687a ) or ( a4678a );
 a4689a <=( a4688a ) or ( a4671a );
 a4690a <=( a4689a ) or ( a4654a );
 a4693a <=( a1118a ) or ( a1119a );
 a4696a <=( a1116a ) or ( a1117a );
 a4697a <=( a4696a ) or ( a4693a );
 a4700a <=( a1114a ) or ( a1115a );
 a4704a <=( a1111a ) or ( a1112a );
 a4705a <=( a1113a ) or ( a4704a );
 a4706a <=( a4705a ) or ( a4700a );
 a4707a <=( a4706a ) or ( a4697a );
 a4710a <=( a1109a ) or ( a1110a );
 a4713a <=( a1107a ) or ( a1108a );
 a4714a <=( a4713a ) or ( a4710a );
 a4717a <=( a1105a ) or ( a1106a );
 a4721a <=( a1102a ) or ( a1103a );
 a4722a <=( a1104a ) or ( a4721a );
 a4723a <=( a4722a ) or ( a4717a );
 a4724a <=( a4723a ) or ( a4714a );
 a4725a <=( a4724a ) or ( a4707a );
 a4728a <=( a1100a ) or ( a1101a );
 a4731a <=( a1098a ) or ( a1099a );
 a4732a <=( a4731a ) or ( a4728a );
 a4735a <=( a1096a ) or ( a1097a );
 a4739a <=( a1093a ) or ( a1094a );
 a4740a <=( a1095a ) or ( a4739a );
 a4741a <=( a4740a ) or ( a4735a );
 a4742a <=( a4741a ) or ( a4732a );
 a4745a <=( a1091a ) or ( a1092a );
 a4748a <=( a1089a ) or ( a1090a );
 a4749a <=( a4748a ) or ( a4745a );
 a4752a <=( a1087a ) or ( a1088a );
 a4756a <=( a1084a ) or ( a1085a );
 a4757a <=( a1086a ) or ( a4756a );
 a4758a <=( a4757a ) or ( a4752a );
 a4759a <=( a4758a ) or ( a4749a );
 a4760a <=( a4759a ) or ( a4742a );
 a4761a <=( a4760a ) or ( a4725a );
 a4762a <=( a4761a ) or ( a4690a );
 a4765a <=( a1082a ) or ( a1083a );
 a4768a <=( a1080a ) or ( a1081a );
 a4769a <=( a4768a ) or ( a4765a );
 a4772a <=( a1078a ) or ( a1079a );
 a4776a <=( a1075a ) or ( a1076a );
 a4777a <=( a1077a ) or ( a4776a );
 a4778a <=( a4777a ) or ( a4772a );
 a4779a <=( a4778a ) or ( a4769a );
 a4782a <=( a1073a ) or ( a1074a );
 a4785a <=( a1071a ) or ( a1072a );
 a4786a <=( a4785a ) or ( a4782a );
 a4789a <=( a1069a ) or ( a1070a );
 a4793a <=( a1066a ) or ( a1067a );
 a4794a <=( a1068a ) or ( a4793a );
 a4795a <=( a4794a ) or ( a4789a );
 a4796a <=( a4795a ) or ( a4786a );
 a4797a <=( a4796a ) or ( a4779a );
 a4800a <=( a1064a ) or ( a1065a );
 a4803a <=( a1062a ) or ( a1063a );
 a4804a <=( a4803a ) or ( a4800a );
 a4807a <=( a1060a ) or ( a1061a );
 a4811a <=( a1057a ) or ( a1058a );
 a4812a <=( a1059a ) or ( a4811a );
 a4813a <=( a4812a ) or ( a4807a );
 a4814a <=( a4813a ) or ( a4804a );
 a4817a <=( a1055a ) or ( a1056a );
 a4820a <=( a1053a ) or ( a1054a );
 a4821a <=( a4820a ) or ( a4817a );
 a4824a <=( a1051a ) or ( a1052a );
 a4828a <=( a1048a ) or ( a1049a );
 a4829a <=( a1050a ) or ( a4828a );
 a4830a <=( a4829a ) or ( a4824a );
 a4831a <=( a4830a ) or ( a4821a );
 a4832a <=( a4831a ) or ( a4814a );
 a4833a <=( a4832a ) or ( a4797a );
 a4836a <=( a1046a ) or ( a1047a );
 a4839a <=( a1044a ) or ( a1045a );
 a4840a <=( a4839a ) or ( a4836a );
 a4843a <=( a1042a ) or ( a1043a );
 a4847a <=( a1039a ) or ( a1040a );
 a4848a <=( a1041a ) or ( a4847a );
 a4849a <=( a4848a ) or ( a4843a );
 a4850a <=( a4849a ) or ( a4840a );
 a4853a <=( a1037a ) or ( a1038a );
 a4856a <=( a1035a ) or ( a1036a );
 a4857a <=( a4856a ) or ( a4853a );
 a4860a <=( a1033a ) or ( a1034a );
 a4864a <=( a1030a ) or ( a1031a );
 a4865a <=( a1032a ) or ( a4864a );
 a4866a <=( a4865a ) or ( a4860a );
 a4867a <=( a4866a ) or ( a4857a );
 a4868a <=( a4867a ) or ( a4850a );
 a4871a <=( a1028a ) or ( a1029a );
 a4874a <=( a1026a ) or ( a1027a );
 a4875a <=( a4874a ) or ( a4871a );
 a4878a <=( a1024a ) or ( a1025a );
 a4882a <=( a1021a ) or ( a1022a );
 a4883a <=( a1023a ) or ( a4882a );
 a4884a <=( a4883a ) or ( a4878a );
 a4885a <=( a4884a ) or ( a4875a );
 a4888a <=( a1019a ) or ( a1020a );
 a4891a <=( a1017a ) or ( a1018a );
 a4892a <=( a4891a ) or ( a4888a );
 a4895a <=( a1015a ) or ( a1016a );
 a4899a <=( a1012a ) or ( a1013a );
 a4900a <=( a1014a ) or ( a4899a );
 a4901a <=( a4900a ) or ( a4895a );
 a4902a <=( a4901a ) or ( a4892a );
 a4903a <=( a4902a ) or ( a4885a );
 a4904a <=( a4903a ) or ( a4868a );
 a4905a <=( a4904a ) or ( a4833a );
 a4906a <=( a4905a ) or ( a4762a );
 a4909a <=( a1010a ) or ( a1011a );
 a4912a <=( a1008a ) or ( a1009a );
 a4913a <=( a4912a ) or ( a4909a );
 a4916a <=( a1006a ) or ( a1007a );
 a4920a <=( a1003a ) or ( a1004a );
 a4921a <=( a1005a ) or ( a4920a );
 a4922a <=( a4921a ) or ( a4916a );
 a4923a <=( a4922a ) or ( a4913a );
 a4926a <=( a1001a ) or ( a1002a );
 a4929a <=( a999a ) or ( a1000a );
 a4930a <=( a4929a ) or ( a4926a );
 a4933a <=( a997a ) or ( a998a );
 a4937a <=( a994a ) or ( a995a );
 a4938a <=( a996a ) or ( a4937a );
 a4939a <=( a4938a ) or ( a4933a );
 a4940a <=( a4939a ) or ( a4930a );
 a4941a <=( a4940a ) or ( a4923a );
 a4944a <=( a992a ) or ( a993a );
 a4947a <=( a990a ) or ( a991a );
 a4948a <=( a4947a ) or ( a4944a );
 a4951a <=( a988a ) or ( a989a );
 a4955a <=( a985a ) or ( a986a );
 a4956a <=( a987a ) or ( a4955a );
 a4957a <=( a4956a ) or ( a4951a );
 a4958a <=( a4957a ) or ( a4948a );
 a4961a <=( a983a ) or ( a984a );
 a4964a <=( a981a ) or ( a982a );
 a4965a <=( a4964a ) or ( a4961a );
 a4968a <=( a979a ) or ( a980a );
 a4972a <=( a976a ) or ( a977a );
 a4973a <=( a978a ) or ( a4972a );
 a4974a <=( a4973a ) or ( a4968a );
 a4975a <=( a4974a ) or ( a4965a );
 a4976a <=( a4975a ) or ( a4958a );
 a4977a <=( a4976a ) or ( a4941a );
 a4980a <=( a974a ) or ( a975a );
 a4983a <=( a972a ) or ( a973a );
 a4984a <=( a4983a ) or ( a4980a );
 a4987a <=( a970a ) or ( a971a );
 a4991a <=( a967a ) or ( a968a );
 a4992a <=( a969a ) or ( a4991a );
 a4993a <=( a4992a ) or ( a4987a );
 a4994a <=( a4993a ) or ( a4984a );
 a4997a <=( a965a ) or ( a966a );
 a5000a <=( a963a ) or ( a964a );
 a5001a <=( a5000a ) or ( a4997a );
 a5004a <=( a961a ) or ( a962a );
 a5008a <=( a958a ) or ( a959a );
 a5009a <=( a960a ) or ( a5008a );
 a5010a <=( a5009a ) or ( a5004a );
 a5011a <=( a5010a ) or ( a5001a );
 a5012a <=( a5011a ) or ( a4994a );
 a5015a <=( a956a ) or ( a957a );
 a5018a <=( a954a ) or ( a955a );
 a5019a <=( a5018a ) or ( a5015a );
 a5022a <=( a952a ) or ( a953a );
 a5026a <=( a949a ) or ( a950a );
 a5027a <=( a951a ) or ( a5026a );
 a5028a <=( a5027a ) or ( a5022a );
 a5029a <=( a5028a ) or ( a5019a );
 a5032a <=( a947a ) or ( a948a );
 a5035a <=( a945a ) or ( a946a );
 a5036a <=( a5035a ) or ( a5032a );
 a5039a <=( a943a ) or ( a944a );
 a5043a <=( a940a ) or ( a941a );
 a5044a <=( a942a ) or ( a5043a );
 a5045a <=( a5044a ) or ( a5039a );
 a5046a <=( a5045a ) or ( a5036a );
 a5047a <=( a5046a ) or ( a5029a );
 a5048a <=( a5047a ) or ( a5012a );
 a5049a <=( a5048a ) or ( a4977a );
 a5052a <=( a938a ) or ( a939a );
 a5055a <=( a936a ) or ( a937a );
 a5056a <=( a5055a ) or ( a5052a );
 a5059a <=( a934a ) or ( a935a );
 a5063a <=( a931a ) or ( a932a );
 a5064a <=( a933a ) or ( a5063a );
 a5065a <=( a5064a ) or ( a5059a );
 a5066a <=( a5065a ) or ( a5056a );
 a5069a <=( a929a ) or ( a930a );
 a5072a <=( a927a ) or ( a928a );
 a5073a <=( a5072a ) or ( a5069a );
 a5076a <=( a925a ) or ( a926a );
 a5080a <=( a922a ) or ( a923a );
 a5081a <=( a924a ) or ( a5080a );
 a5082a <=( a5081a ) or ( a5076a );
 a5083a <=( a5082a ) or ( a5073a );
 a5084a <=( a5083a ) or ( a5066a );
 a5087a <=( a920a ) or ( a921a );
 a5090a <=( a918a ) or ( a919a );
 a5091a <=( a5090a ) or ( a5087a );
 a5094a <=( a916a ) or ( a917a );
 a5098a <=( a913a ) or ( a914a );
 a5099a <=( a915a ) or ( a5098a );
 a5100a <=( a5099a ) or ( a5094a );
 a5101a <=( a5100a ) or ( a5091a );
 a5104a <=( a911a ) or ( a912a );
 a5107a <=( a909a ) or ( a910a );
 a5108a <=( a5107a ) or ( a5104a );
 a5111a <=( a907a ) or ( a908a );
 a5115a <=( a904a ) or ( a905a );
 a5116a <=( a906a ) or ( a5115a );
 a5117a <=( a5116a ) or ( a5111a );
 a5118a <=( a5117a ) or ( a5108a );
 a5119a <=( a5118a ) or ( a5101a );
 a5120a <=( a5119a ) or ( a5084a );
 a5123a <=( a902a ) or ( a903a );
 a5126a <=( a900a ) or ( a901a );
 a5127a <=( a5126a ) or ( a5123a );
 a5130a <=( a898a ) or ( a899a );
 a5134a <=( a895a ) or ( a896a );
 a5135a <=( a897a ) or ( a5134a );
 a5136a <=( a5135a ) or ( a5130a );
 a5137a <=( a5136a ) or ( a5127a );
 a5140a <=( a893a ) or ( a894a );
 a5143a <=( a891a ) or ( a892a );
 a5144a <=( a5143a ) or ( a5140a );
 a5147a <=( a889a ) or ( a890a );
 a5151a <=( a886a ) or ( a887a );
 a5152a <=( a888a ) or ( a5151a );
 a5153a <=( a5152a ) or ( a5147a );
 a5154a <=( a5153a ) or ( a5144a );
 a5155a <=( a5154a ) or ( a5137a );
 a5158a <=( a884a ) or ( a885a );
 a5161a <=( a882a ) or ( a883a );
 a5162a <=( a5161a ) or ( a5158a );
 a5165a <=( a880a ) or ( a881a );
 a5169a <=( a877a ) or ( a878a );
 a5170a <=( a879a ) or ( a5169a );
 a5171a <=( a5170a ) or ( a5165a );
 a5172a <=( a5171a ) or ( a5162a );
 a5175a <=( a875a ) or ( a876a );
 a5178a <=( a873a ) or ( a874a );
 a5179a <=( a5178a ) or ( a5175a );
 a5182a <=( a871a ) or ( a872a );
 a5186a <=( a868a ) or ( a869a );
 a5187a <=( a870a ) or ( a5186a );
 a5188a <=( a5187a ) or ( a5182a );
 a5189a <=( a5188a ) or ( a5179a );
 a5190a <=( a5189a ) or ( a5172a );
 a5191a <=( a5190a ) or ( a5155a );
 a5192a <=( a5191a ) or ( a5120a );
 a5193a <=( a5192a ) or ( a5049a );
 a5194a <=( a5193a ) or ( a4906a );
 a5197a <=( a866a ) or ( a867a );
 a5200a <=( a864a ) or ( a865a );
 a5201a <=( a5200a ) or ( a5197a );
 a5204a <=( a862a ) or ( a863a );
 a5208a <=( a859a ) or ( a860a );
 a5209a <=( a861a ) or ( a5208a );
 a5210a <=( a5209a ) or ( a5204a );
 a5211a <=( a5210a ) or ( a5201a );
 a5214a <=( a857a ) or ( a858a );
 a5217a <=( a855a ) or ( a856a );
 a5218a <=( a5217a ) or ( a5214a );
 a5221a <=( a853a ) or ( a854a );
 a5225a <=( a850a ) or ( a851a );
 a5226a <=( a852a ) or ( a5225a );
 a5227a <=( a5226a ) or ( a5221a );
 a5228a <=( a5227a ) or ( a5218a );
 a5229a <=( a5228a ) or ( a5211a );
 a5232a <=( a848a ) or ( a849a );
 a5235a <=( a846a ) or ( a847a );
 a5236a <=( a5235a ) or ( a5232a );
 a5239a <=( a844a ) or ( a845a );
 a5243a <=( a841a ) or ( a842a );
 a5244a <=( a843a ) or ( a5243a );
 a5245a <=( a5244a ) or ( a5239a );
 a5246a <=( a5245a ) or ( a5236a );
 a5249a <=( a839a ) or ( a840a );
 a5252a <=( a837a ) or ( a838a );
 a5253a <=( a5252a ) or ( a5249a );
 a5256a <=( a835a ) or ( a836a );
 a5260a <=( a832a ) or ( a833a );
 a5261a <=( a834a ) or ( a5260a );
 a5262a <=( a5261a ) or ( a5256a );
 a5263a <=( a5262a ) or ( a5253a );
 a5264a <=( a5263a ) or ( a5246a );
 a5265a <=( a5264a ) or ( a5229a );
 a5268a <=( a830a ) or ( a831a );
 a5271a <=( a828a ) or ( a829a );
 a5272a <=( a5271a ) or ( a5268a );
 a5275a <=( a826a ) or ( a827a );
 a5279a <=( a823a ) or ( a824a );
 a5280a <=( a825a ) or ( a5279a );
 a5281a <=( a5280a ) or ( a5275a );
 a5282a <=( a5281a ) or ( a5272a );
 a5285a <=( a821a ) or ( a822a );
 a5288a <=( a819a ) or ( a820a );
 a5289a <=( a5288a ) or ( a5285a );
 a5292a <=( a817a ) or ( a818a );
 a5296a <=( a814a ) or ( a815a );
 a5297a <=( a816a ) or ( a5296a );
 a5298a <=( a5297a ) or ( a5292a );
 a5299a <=( a5298a ) or ( a5289a );
 a5300a <=( a5299a ) or ( a5282a );
 a5303a <=( a812a ) or ( a813a );
 a5306a <=( a810a ) or ( a811a );
 a5307a <=( a5306a ) or ( a5303a );
 a5310a <=( a808a ) or ( a809a );
 a5314a <=( a805a ) or ( a806a );
 a5315a <=( a807a ) or ( a5314a );
 a5316a <=( a5315a ) or ( a5310a );
 a5317a <=( a5316a ) or ( a5307a );
 a5320a <=( a803a ) or ( a804a );
 a5323a <=( a801a ) or ( a802a );
 a5324a <=( a5323a ) or ( a5320a );
 a5327a <=( a799a ) or ( a800a );
 a5331a <=( a796a ) or ( a797a );
 a5332a <=( a798a ) or ( a5331a );
 a5333a <=( a5332a ) or ( a5327a );
 a5334a <=( a5333a ) or ( a5324a );
 a5335a <=( a5334a ) or ( a5317a );
 a5336a <=( a5335a ) or ( a5300a );
 a5337a <=( a5336a ) or ( a5265a );
 a5340a <=( a794a ) or ( a795a );
 a5343a <=( a792a ) or ( a793a );
 a5344a <=( a5343a ) or ( a5340a );
 a5347a <=( a790a ) or ( a791a );
 a5351a <=( a787a ) or ( a788a );
 a5352a <=( a789a ) or ( a5351a );
 a5353a <=( a5352a ) or ( a5347a );
 a5354a <=( a5353a ) or ( a5344a );
 a5357a <=( a785a ) or ( a786a );
 a5360a <=( a783a ) or ( a784a );
 a5361a <=( a5360a ) or ( a5357a );
 a5364a <=( a781a ) or ( a782a );
 a5368a <=( a778a ) or ( a779a );
 a5369a <=( a780a ) or ( a5368a );
 a5370a <=( a5369a ) or ( a5364a );
 a5371a <=( a5370a ) or ( a5361a );
 a5372a <=( a5371a ) or ( a5354a );
 a5375a <=( a776a ) or ( a777a );
 a5378a <=( a774a ) or ( a775a );
 a5379a <=( a5378a ) or ( a5375a );
 a5382a <=( a772a ) or ( a773a );
 a5386a <=( a769a ) or ( a770a );
 a5387a <=( a771a ) or ( a5386a );
 a5388a <=( a5387a ) or ( a5382a );
 a5389a <=( a5388a ) or ( a5379a );
 a5392a <=( a767a ) or ( a768a );
 a5395a <=( a765a ) or ( a766a );
 a5396a <=( a5395a ) or ( a5392a );
 a5399a <=( a763a ) or ( a764a );
 a5403a <=( a760a ) or ( a761a );
 a5404a <=( a762a ) or ( a5403a );
 a5405a <=( a5404a ) or ( a5399a );
 a5406a <=( a5405a ) or ( a5396a );
 a5407a <=( a5406a ) or ( a5389a );
 a5408a <=( a5407a ) or ( a5372a );
 a5411a <=( a758a ) or ( a759a );
 a5414a <=( a756a ) or ( a757a );
 a5415a <=( a5414a ) or ( a5411a );
 a5418a <=( a754a ) or ( a755a );
 a5422a <=( a751a ) or ( a752a );
 a5423a <=( a753a ) or ( a5422a );
 a5424a <=( a5423a ) or ( a5418a );
 a5425a <=( a5424a ) or ( a5415a );
 a5428a <=( a749a ) or ( a750a );
 a5431a <=( a747a ) or ( a748a );
 a5432a <=( a5431a ) or ( a5428a );
 a5435a <=( a745a ) or ( a746a );
 a5439a <=( a742a ) or ( a743a );
 a5440a <=( a744a ) or ( a5439a );
 a5441a <=( a5440a ) or ( a5435a );
 a5442a <=( a5441a ) or ( a5432a );
 a5443a <=( a5442a ) or ( a5425a );
 a5446a <=( a740a ) or ( a741a );
 a5449a <=( a738a ) or ( a739a );
 a5450a <=( a5449a ) or ( a5446a );
 a5453a <=( a736a ) or ( a737a );
 a5457a <=( a733a ) or ( a734a );
 a5458a <=( a735a ) or ( a5457a );
 a5459a <=( a5458a ) or ( a5453a );
 a5460a <=( a5459a ) or ( a5450a );
 a5463a <=( a731a ) or ( a732a );
 a5466a <=( a729a ) or ( a730a );
 a5467a <=( a5466a ) or ( a5463a );
 a5470a <=( a727a ) or ( a728a );
 a5474a <=( a724a ) or ( a725a );
 a5475a <=( a726a ) or ( a5474a );
 a5476a <=( a5475a ) or ( a5470a );
 a5477a <=( a5476a ) or ( a5467a );
 a5478a <=( a5477a ) or ( a5460a );
 a5479a <=( a5478a ) or ( a5443a );
 a5480a <=( a5479a ) or ( a5408a );
 a5481a <=( a5480a ) or ( a5337a );
 a5484a <=( a722a ) or ( a723a );
 a5487a <=( a720a ) or ( a721a );
 a5488a <=( a5487a ) or ( a5484a );
 a5491a <=( a718a ) or ( a719a );
 a5495a <=( a715a ) or ( a716a );
 a5496a <=( a717a ) or ( a5495a );
 a5497a <=( a5496a ) or ( a5491a );
 a5498a <=( a5497a ) or ( a5488a );
 a5501a <=( a713a ) or ( a714a );
 a5504a <=( a711a ) or ( a712a );
 a5505a <=( a5504a ) or ( a5501a );
 a5508a <=( a709a ) or ( a710a );
 a5512a <=( a706a ) or ( a707a );
 a5513a <=( a708a ) or ( a5512a );
 a5514a <=( a5513a ) or ( a5508a );
 a5515a <=( a5514a ) or ( a5505a );
 a5516a <=( a5515a ) or ( a5498a );
 a5519a <=( a704a ) or ( a705a );
 a5522a <=( a702a ) or ( a703a );
 a5523a <=( a5522a ) or ( a5519a );
 a5526a <=( a700a ) or ( a701a );
 a5530a <=( a697a ) or ( a698a );
 a5531a <=( a699a ) or ( a5530a );
 a5532a <=( a5531a ) or ( a5526a );
 a5533a <=( a5532a ) or ( a5523a );
 a5536a <=( a695a ) or ( a696a );
 a5539a <=( a693a ) or ( a694a );
 a5540a <=( a5539a ) or ( a5536a );
 a5543a <=( a691a ) or ( a692a );
 a5547a <=( a688a ) or ( a689a );
 a5548a <=( a690a ) or ( a5547a );
 a5549a <=( a5548a ) or ( a5543a );
 a5550a <=( a5549a ) or ( a5540a );
 a5551a <=( a5550a ) or ( a5533a );
 a5552a <=( a5551a ) or ( a5516a );
 a5555a <=( a686a ) or ( a687a );
 a5558a <=( a684a ) or ( a685a );
 a5559a <=( a5558a ) or ( a5555a );
 a5562a <=( a682a ) or ( a683a );
 a5566a <=( a679a ) or ( a680a );
 a5567a <=( a681a ) or ( a5566a );
 a5568a <=( a5567a ) or ( a5562a );
 a5569a <=( a5568a ) or ( a5559a );
 a5572a <=( a677a ) or ( a678a );
 a5575a <=( a675a ) or ( a676a );
 a5576a <=( a5575a ) or ( a5572a );
 a5579a <=( a673a ) or ( a674a );
 a5583a <=( a670a ) or ( a671a );
 a5584a <=( a672a ) or ( a5583a );
 a5585a <=( a5584a ) or ( a5579a );
 a5586a <=( a5585a ) or ( a5576a );
 a5587a <=( a5586a ) or ( a5569a );
 a5590a <=( a668a ) or ( a669a );
 a5593a <=( a666a ) or ( a667a );
 a5594a <=( a5593a ) or ( a5590a );
 a5597a <=( a664a ) or ( a665a );
 a5601a <=( a661a ) or ( a662a );
 a5602a <=( a663a ) or ( a5601a );
 a5603a <=( a5602a ) or ( a5597a );
 a5604a <=( a5603a ) or ( a5594a );
 a5607a <=( a659a ) or ( a660a );
 a5610a <=( a657a ) or ( a658a );
 a5611a <=( a5610a ) or ( a5607a );
 a5614a <=( a655a ) or ( a656a );
 a5618a <=( a652a ) or ( a653a );
 a5619a <=( a654a ) or ( a5618a );
 a5620a <=( a5619a ) or ( a5614a );
 a5621a <=( a5620a ) or ( a5611a );
 a5622a <=( a5621a ) or ( a5604a );
 a5623a <=( a5622a ) or ( a5587a );
 a5624a <=( a5623a ) or ( a5552a );
 a5627a <=( a650a ) or ( a651a );
 a5630a <=( a648a ) or ( a649a );
 a5631a <=( a5630a ) or ( a5627a );
 a5634a <=( a646a ) or ( a647a );
 a5638a <=( a643a ) or ( a644a );
 a5639a <=( a645a ) or ( a5638a );
 a5640a <=( a5639a ) or ( a5634a );
 a5641a <=( a5640a ) or ( a5631a );
 a5644a <=( a641a ) or ( a642a );
 a5647a <=( a639a ) or ( a640a );
 a5648a <=( a5647a ) or ( a5644a );
 a5651a <=( a637a ) or ( a638a );
 a5655a <=( a634a ) or ( a635a );
 a5656a <=( a636a ) or ( a5655a );
 a5657a <=( a5656a ) or ( a5651a );
 a5658a <=( a5657a ) or ( a5648a );
 a5659a <=( a5658a ) or ( a5641a );
 a5662a <=( a632a ) or ( a633a );
 a5665a <=( a630a ) or ( a631a );
 a5666a <=( a5665a ) or ( a5662a );
 a5669a <=( a628a ) or ( a629a );
 a5673a <=( a625a ) or ( a626a );
 a5674a <=( a627a ) or ( a5673a );
 a5675a <=( a5674a ) or ( a5669a );
 a5676a <=( a5675a ) or ( a5666a );
 a5679a <=( a623a ) or ( a624a );
 a5682a <=( a621a ) or ( a622a );
 a5683a <=( a5682a ) or ( a5679a );
 a5686a <=( a619a ) or ( a620a );
 a5690a <=( a616a ) or ( a617a );
 a5691a <=( a618a ) or ( a5690a );
 a5692a <=( a5691a ) or ( a5686a );
 a5693a <=( a5692a ) or ( a5683a );
 a5694a <=( a5693a ) or ( a5676a );
 a5695a <=( a5694a ) or ( a5659a );
 a5698a <=( a614a ) or ( a615a );
 a5701a <=( a612a ) or ( a613a );
 a5702a <=( a5701a ) or ( a5698a );
 a5705a <=( a610a ) or ( a611a );
 a5709a <=( a607a ) or ( a608a );
 a5710a <=( a609a ) or ( a5709a );
 a5711a <=( a5710a ) or ( a5705a );
 a5712a <=( a5711a ) or ( a5702a );
 a5715a <=( a605a ) or ( a606a );
 a5718a <=( a603a ) or ( a604a );
 a5719a <=( a5718a ) or ( a5715a );
 a5722a <=( a601a ) or ( a602a );
 a5726a <=( a598a ) or ( a599a );
 a5727a <=( a600a ) or ( a5726a );
 a5728a <=( a5727a ) or ( a5722a );
 a5729a <=( a5728a ) or ( a5719a );
 a5730a <=( a5729a ) or ( a5712a );
 a5733a <=( a596a ) or ( a597a );
 a5736a <=( a594a ) or ( a595a );
 a5737a <=( a5736a ) or ( a5733a );
 a5740a <=( a592a ) or ( a593a );
 a5744a <=( a589a ) or ( a590a );
 a5745a <=( a591a ) or ( a5744a );
 a5746a <=( a5745a ) or ( a5740a );
 a5747a <=( a5746a ) or ( a5737a );
 a5750a <=( a587a ) or ( a588a );
 a5754a <=( a584a ) or ( a585a );
 a5755a <=( a586a ) or ( a5754a );
 a5756a <=( a5755a ) or ( a5750a );
 a5759a <=( a582a ) or ( a583a );
 a5763a <=( a579a ) or ( a580a );
 a5764a <=( a581a ) or ( a5763a );
 a5765a <=( a5764a ) or ( a5759a );
 a5766a <=( a5765a ) or ( a5756a );
 a5767a <=( a5766a ) or ( a5747a );
 a5768a <=( a5767a ) or ( a5730a );
 a5769a <=( a5768a ) or ( a5695a );
 a5770a <=( a5769a ) or ( a5624a );
 a5771a <=( a5770a ) or ( a5481a );
 a5772a <=( a5771a ) or ( a5194a );
 a5775a <=( a577a ) or ( a578a );
 a5778a <=( a575a ) or ( a576a );
 a5779a <=( a5778a ) or ( a5775a );
 a5782a <=( a573a ) or ( a574a );
 a5786a <=( a570a ) or ( a571a );
 a5787a <=( a572a ) or ( a5786a );
 a5788a <=( a5787a ) or ( a5782a );
 a5789a <=( a5788a ) or ( a5779a );
 a5792a <=( a568a ) or ( a569a );
 a5795a <=( a566a ) or ( a567a );
 a5796a <=( a5795a ) or ( a5792a );
 a5799a <=( a564a ) or ( a565a );
 a5803a <=( a561a ) or ( a562a );
 a5804a <=( a563a ) or ( a5803a );
 a5805a <=( a5804a ) or ( a5799a );
 a5806a <=( a5805a ) or ( a5796a );
 a5807a <=( a5806a ) or ( a5789a );
 a5810a <=( a559a ) or ( a560a );
 a5813a <=( a557a ) or ( a558a );
 a5814a <=( a5813a ) or ( a5810a );
 a5817a <=( a555a ) or ( a556a );
 a5821a <=( a552a ) or ( a553a );
 a5822a <=( a554a ) or ( a5821a );
 a5823a <=( a5822a ) or ( a5817a );
 a5824a <=( a5823a ) or ( a5814a );
 a5827a <=( a550a ) or ( a551a );
 a5830a <=( a548a ) or ( a549a );
 a5831a <=( a5830a ) or ( a5827a );
 a5834a <=( a546a ) or ( a547a );
 a5838a <=( a543a ) or ( a544a );
 a5839a <=( a545a ) or ( a5838a );
 a5840a <=( a5839a ) or ( a5834a );
 a5841a <=( a5840a ) or ( a5831a );
 a5842a <=( a5841a ) or ( a5824a );
 a5843a <=( a5842a ) or ( a5807a );
 a5846a <=( a541a ) or ( a542a );
 a5849a <=( a539a ) or ( a540a );
 a5850a <=( a5849a ) or ( a5846a );
 a5853a <=( a537a ) or ( a538a );
 a5857a <=( a534a ) or ( a535a );
 a5858a <=( a536a ) or ( a5857a );
 a5859a <=( a5858a ) or ( a5853a );
 a5860a <=( a5859a ) or ( a5850a );
 a5863a <=( a532a ) or ( a533a );
 a5866a <=( a530a ) or ( a531a );
 a5867a <=( a5866a ) or ( a5863a );
 a5870a <=( a528a ) or ( a529a );
 a5874a <=( a525a ) or ( a526a );
 a5875a <=( a527a ) or ( a5874a );
 a5876a <=( a5875a ) or ( a5870a );
 a5877a <=( a5876a ) or ( a5867a );
 a5878a <=( a5877a ) or ( a5860a );
 a5881a <=( a523a ) or ( a524a );
 a5884a <=( a521a ) or ( a522a );
 a5885a <=( a5884a ) or ( a5881a );
 a5888a <=( a519a ) or ( a520a );
 a5892a <=( a516a ) or ( a517a );
 a5893a <=( a518a ) or ( a5892a );
 a5894a <=( a5893a ) or ( a5888a );
 a5895a <=( a5894a ) or ( a5885a );
 a5898a <=( a514a ) or ( a515a );
 a5901a <=( a512a ) or ( a513a );
 a5902a <=( a5901a ) or ( a5898a );
 a5905a <=( a510a ) or ( a511a );
 a5909a <=( a507a ) or ( a508a );
 a5910a <=( a509a ) or ( a5909a );
 a5911a <=( a5910a ) or ( a5905a );
 a5912a <=( a5911a ) or ( a5902a );
 a5913a <=( a5912a ) or ( a5895a );
 a5914a <=( a5913a ) or ( a5878a );
 a5915a <=( a5914a ) or ( a5843a );
 a5918a <=( a505a ) or ( a506a );
 a5921a <=( a503a ) or ( a504a );
 a5922a <=( a5921a ) or ( a5918a );
 a5925a <=( a501a ) or ( a502a );
 a5929a <=( a498a ) or ( a499a );
 a5930a <=( a500a ) or ( a5929a );
 a5931a <=( a5930a ) or ( a5925a );
 a5932a <=( a5931a ) or ( a5922a );
 a5935a <=( a496a ) or ( a497a );
 a5938a <=( a494a ) or ( a495a );
 a5939a <=( a5938a ) or ( a5935a );
 a5942a <=( a492a ) or ( a493a );
 a5946a <=( a489a ) or ( a490a );
 a5947a <=( a491a ) or ( a5946a );
 a5948a <=( a5947a ) or ( a5942a );
 a5949a <=( a5948a ) or ( a5939a );
 a5950a <=( a5949a ) or ( a5932a );
 a5953a <=( a487a ) or ( a488a );
 a5956a <=( a485a ) or ( a486a );
 a5957a <=( a5956a ) or ( a5953a );
 a5960a <=( a483a ) or ( a484a );
 a5964a <=( a480a ) or ( a481a );
 a5965a <=( a482a ) or ( a5964a );
 a5966a <=( a5965a ) or ( a5960a );
 a5967a <=( a5966a ) or ( a5957a );
 a5970a <=( a478a ) or ( a479a );
 a5973a <=( a476a ) or ( a477a );
 a5974a <=( a5973a ) or ( a5970a );
 a5977a <=( a474a ) or ( a475a );
 a5981a <=( a471a ) or ( a472a );
 a5982a <=( a473a ) or ( a5981a );
 a5983a <=( a5982a ) or ( a5977a );
 a5984a <=( a5983a ) or ( a5974a );
 a5985a <=( a5984a ) or ( a5967a );
 a5986a <=( a5985a ) or ( a5950a );
 a5989a <=( a469a ) or ( a470a );
 a5992a <=( a467a ) or ( a468a );
 a5993a <=( a5992a ) or ( a5989a );
 a5996a <=( a465a ) or ( a466a );
 a6000a <=( a462a ) or ( a463a );
 a6001a <=( a464a ) or ( a6000a );
 a6002a <=( a6001a ) or ( a5996a );
 a6003a <=( a6002a ) or ( a5993a );
 a6006a <=( a460a ) or ( a461a );
 a6009a <=( a458a ) or ( a459a );
 a6010a <=( a6009a ) or ( a6006a );
 a6013a <=( a456a ) or ( a457a );
 a6017a <=( a453a ) or ( a454a );
 a6018a <=( a455a ) or ( a6017a );
 a6019a <=( a6018a ) or ( a6013a );
 a6020a <=( a6019a ) or ( a6010a );
 a6021a <=( a6020a ) or ( a6003a );
 a6024a <=( a451a ) or ( a452a );
 a6027a <=( a449a ) or ( a450a );
 a6028a <=( a6027a ) or ( a6024a );
 a6031a <=( a447a ) or ( a448a );
 a6035a <=( a444a ) or ( a445a );
 a6036a <=( a446a ) or ( a6035a );
 a6037a <=( a6036a ) or ( a6031a );
 a6038a <=( a6037a ) or ( a6028a );
 a6041a <=( a442a ) or ( a443a );
 a6044a <=( a440a ) or ( a441a );
 a6045a <=( a6044a ) or ( a6041a );
 a6048a <=( a438a ) or ( a439a );
 a6052a <=( a435a ) or ( a436a );
 a6053a <=( a437a ) or ( a6052a );
 a6054a <=( a6053a ) or ( a6048a );
 a6055a <=( a6054a ) or ( a6045a );
 a6056a <=( a6055a ) or ( a6038a );
 a6057a <=( a6056a ) or ( a6021a );
 a6058a <=( a6057a ) or ( a5986a );
 a6059a <=( a6058a ) or ( a5915a );
 a6062a <=( a433a ) or ( a434a );
 a6065a <=( a431a ) or ( a432a );
 a6066a <=( a6065a ) or ( a6062a );
 a6069a <=( a429a ) or ( a430a );
 a6073a <=( a426a ) or ( a427a );
 a6074a <=( a428a ) or ( a6073a );
 a6075a <=( a6074a ) or ( a6069a );
 a6076a <=( a6075a ) or ( a6066a );
 a6079a <=( a424a ) or ( a425a );
 a6082a <=( a422a ) or ( a423a );
 a6083a <=( a6082a ) or ( a6079a );
 a6086a <=( a420a ) or ( a421a );
 a6090a <=( a417a ) or ( a418a );
 a6091a <=( a419a ) or ( a6090a );
 a6092a <=( a6091a ) or ( a6086a );
 a6093a <=( a6092a ) or ( a6083a );
 a6094a <=( a6093a ) or ( a6076a );
 a6097a <=( a415a ) or ( a416a );
 a6100a <=( a413a ) or ( a414a );
 a6101a <=( a6100a ) or ( a6097a );
 a6104a <=( a411a ) or ( a412a );
 a6108a <=( a408a ) or ( a409a );
 a6109a <=( a410a ) or ( a6108a );
 a6110a <=( a6109a ) or ( a6104a );
 a6111a <=( a6110a ) or ( a6101a );
 a6114a <=( a406a ) or ( a407a );
 a6117a <=( a404a ) or ( a405a );
 a6118a <=( a6117a ) or ( a6114a );
 a6121a <=( a402a ) or ( a403a );
 a6125a <=( a399a ) or ( a400a );
 a6126a <=( a401a ) or ( a6125a );
 a6127a <=( a6126a ) or ( a6121a );
 a6128a <=( a6127a ) or ( a6118a );
 a6129a <=( a6128a ) or ( a6111a );
 a6130a <=( a6129a ) or ( a6094a );
 a6133a <=( a397a ) or ( a398a );
 a6136a <=( a395a ) or ( a396a );
 a6137a <=( a6136a ) or ( a6133a );
 a6140a <=( a393a ) or ( a394a );
 a6144a <=( a390a ) or ( a391a );
 a6145a <=( a392a ) or ( a6144a );
 a6146a <=( a6145a ) or ( a6140a );
 a6147a <=( a6146a ) or ( a6137a );
 a6150a <=( a388a ) or ( a389a );
 a6153a <=( a386a ) or ( a387a );
 a6154a <=( a6153a ) or ( a6150a );
 a6157a <=( a384a ) or ( a385a );
 a6161a <=( a381a ) or ( a382a );
 a6162a <=( a383a ) or ( a6161a );
 a6163a <=( a6162a ) or ( a6157a );
 a6164a <=( a6163a ) or ( a6154a );
 a6165a <=( a6164a ) or ( a6147a );
 a6168a <=( a379a ) or ( a380a );
 a6171a <=( a377a ) or ( a378a );
 a6172a <=( a6171a ) or ( a6168a );
 a6175a <=( a375a ) or ( a376a );
 a6179a <=( a372a ) or ( a373a );
 a6180a <=( a374a ) or ( a6179a );
 a6181a <=( a6180a ) or ( a6175a );
 a6182a <=( a6181a ) or ( a6172a );
 a6185a <=( a370a ) or ( a371a );
 a6188a <=( a368a ) or ( a369a );
 a6189a <=( a6188a ) or ( a6185a );
 a6192a <=( a366a ) or ( a367a );
 a6196a <=( a363a ) or ( a364a );
 a6197a <=( a365a ) or ( a6196a );
 a6198a <=( a6197a ) or ( a6192a );
 a6199a <=( a6198a ) or ( a6189a );
 a6200a <=( a6199a ) or ( a6182a );
 a6201a <=( a6200a ) or ( a6165a );
 a6202a <=( a6201a ) or ( a6130a );
 a6205a <=( a361a ) or ( a362a );
 a6208a <=( a359a ) or ( a360a );
 a6209a <=( a6208a ) or ( a6205a );
 a6212a <=( a357a ) or ( a358a );
 a6216a <=( a354a ) or ( a355a );
 a6217a <=( a356a ) or ( a6216a );
 a6218a <=( a6217a ) or ( a6212a );
 a6219a <=( a6218a ) or ( a6209a );
 a6222a <=( a352a ) or ( a353a );
 a6225a <=( a350a ) or ( a351a );
 a6226a <=( a6225a ) or ( a6222a );
 a6229a <=( a348a ) or ( a349a );
 a6233a <=( a345a ) or ( a346a );
 a6234a <=( a347a ) or ( a6233a );
 a6235a <=( a6234a ) or ( a6229a );
 a6236a <=( a6235a ) or ( a6226a );
 a6237a <=( a6236a ) or ( a6219a );
 a6240a <=( a343a ) or ( a344a );
 a6243a <=( a341a ) or ( a342a );
 a6244a <=( a6243a ) or ( a6240a );
 a6247a <=( a339a ) or ( a340a );
 a6251a <=( a336a ) or ( a337a );
 a6252a <=( a338a ) or ( a6251a );
 a6253a <=( a6252a ) or ( a6247a );
 a6254a <=( a6253a ) or ( a6244a );
 a6257a <=( a334a ) or ( a335a );
 a6260a <=( a332a ) or ( a333a );
 a6261a <=( a6260a ) or ( a6257a );
 a6264a <=( a330a ) or ( a331a );
 a6268a <=( a327a ) or ( a328a );
 a6269a <=( a329a ) or ( a6268a );
 a6270a <=( a6269a ) or ( a6264a );
 a6271a <=( a6270a ) or ( a6261a );
 a6272a <=( a6271a ) or ( a6254a );
 a6273a <=( a6272a ) or ( a6237a );
 a6276a <=( a325a ) or ( a326a );
 a6279a <=( a323a ) or ( a324a );
 a6280a <=( a6279a ) or ( a6276a );
 a6283a <=( a321a ) or ( a322a );
 a6287a <=( a318a ) or ( a319a );
 a6288a <=( a320a ) or ( a6287a );
 a6289a <=( a6288a ) or ( a6283a );
 a6290a <=( a6289a ) or ( a6280a );
 a6293a <=( a316a ) or ( a317a );
 a6296a <=( a314a ) or ( a315a );
 a6297a <=( a6296a ) or ( a6293a );
 a6300a <=( a312a ) or ( a313a );
 a6304a <=( a309a ) or ( a310a );
 a6305a <=( a311a ) or ( a6304a );
 a6306a <=( a6305a ) or ( a6300a );
 a6307a <=( a6306a ) or ( a6297a );
 a6308a <=( a6307a ) or ( a6290a );
 a6311a <=( a307a ) or ( a308a );
 a6314a <=( a305a ) or ( a306a );
 a6315a <=( a6314a ) or ( a6311a );
 a6318a <=( a303a ) or ( a304a );
 a6322a <=( a300a ) or ( a301a );
 a6323a <=( a302a ) or ( a6322a );
 a6324a <=( a6323a ) or ( a6318a );
 a6325a <=( a6324a ) or ( a6315a );
 a6328a <=( a298a ) or ( a299a );
 a6332a <=( a295a ) or ( a296a );
 a6333a <=( a297a ) or ( a6332a );
 a6334a <=( a6333a ) or ( a6328a );
 a6337a <=( a293a ) or ( a294a );
 a6341a <=( a290a ) or ( a291a );
 a6342a <=( a292a ) or ( a6341a );
 a6343a <=( a6342a ) or ( a6337a );
 a6344a <=( a6343a ) or ( a6334a );
 a6345a <=( a6344a ) or ( a6325a );
 a6346a <=( a6345a ) or ( a6308a );
 a6347a <=( a6346a ) or ( a6273a );
 a6348a <=( a6347a ) or ( a6202a );
 a6349a <=( a6348a ) or ( a6059a );
 a6352a <=( a288a ) or ( a289a );
 a6355a <=( a286a ) or ( a287a );
 a6356a <=( a6355a ) or ( a6352a );
 a6359a <=( a284a ) or ( a285a );
 a6363a <=( a281a ) or ( a282a );
 a6364a <=( a283a ) or ( a6363a );
 a6365a <=( a6364a ) or ( a6359a );
 a6366a <=( a6365a ) or ( a6356a );
 a6369a <=( a279a ) or ( a280a );
 a6372a <=( a277a ) or ( a278a );
 a6373a <=( a6372a ) or ( a6369a );
 a6376a <=( a275a ) or ( a276a );
 a6380a <=( a272a ) or ( a273a );
 a6381a <=( a274a ) or ( a6380a );
 a6382a <=( a6381a ) or ( a6376a );
 a6383a <=( a6382a ) or ( a6373a );
 a6384a <=( a6383a ) or ( a6366a );
 a6387a <=( a270a ) or ( a271a );
 a6390a <=( a268a ) or ( a269a );
 a6391a <=( a6390a ) or ( a6387a );
 a6394a <=( a266a ) or ( a267a );
 a6398a <=( a263a ) or ( a264a );
 a6399a <=( a265a ) or ( a6398a );
 a6400a <=( a6399a ) or ( a6394a );
 a6401a <=( a6400a ) or ( a6391a );
 a6404a <=( a261a ) or ( a262a );
 a6407a <=( a259a ) or ( a260a );
 a6408a <=( a6407a ) or ( a6404a );
 a6411a <=( a257a ) or ( a258a );
 a6415a <=( a254a ) or ( a255a );
 a6416a <=( a256a ) or ( a6415a );
 a6417a <=( a6416a ) or ( a6411a );
 a6418a <=( a6417a ) or ( a6408a );
 a6419a <=( a6418a ) or ( a6401a );
 a6420a <=( a6419a ) or ( a6384a );
 a6423a <=( a252a ) or ( a253a );
 a6426a <=( a250a ) or ( a251a );
 a6427a <=( a6426a ) or ( a6423a );
 a6430a <=( a248a ) or ( a249a );
 a6434a <=( a245a ) or ( a246a );
 a6435a <=( a247a ) or ( a6434a );
 a6436a <=( a6435a ) or ( a6430a );
 a6437a <=( a6436a ) or ( a6427a );
 a6440a <=( a243a ) or ( a244a );
 a6443a <=( a241a ) or ( a242a );
 a6444a <=( a6443a ) or ( a6440a );
 a6447a <=( a239a ) or ( a240a );
 a6451a <=( a236a ) or ( a237a );
 a6452a <=( a238a ) or ( a6451a );
 a6453a <=( a6452a ) or ( a6447a );
 a6454a <=( a6453a ) or ( a6444a );
 a6455a <=( a6454a ) or ( a6437a );
 a6458a <=( a234a ) or ( a235a );
 a6461a <=( a232a ) or ( a233a );
 a6462a <=( a6461a ) or ( a6458a );
 a6465a <=( a230a ) or ( a231a );
 a6469a <=( a227a ) or ( a228a );
 a6470a <=( a229a ) or ( a6469a );
 a6471a <=( a6470a ) or ( a6465a );
 a6472a <=( a6471a ) or ( a6462a );
 a6475a <=( a225a ) or ( a226a );
 a6478a <=( a223a ) or ( a224a );
 a6479a <=( a6478a ) or ( a6475a );
 a6482a <=( a221a ) or ( a222a );
 a6486a <=( a218a ) or ( a219a );
 a6487a <=( a220a ) or ( a6486a );
 a6488a <=( a6487a ) or ( a6482a );
 a6489a <=( a6488a ) or ( a6479a );
 a6490a <=( a6489a ) or ( a6472a );
 a6491a <=( a6490a ) or ( a6455a );
 a6492a <=( a6491a ) or ( a6420a );
 a6495a <=( a216a ) or ( a217a );
 a6498a <=( a214a ) or ( a215a );
 a6499a <=( a6498a ) or ( a6495a );
 a6502a <=( a212a ) or ( a213a );
 a6506a <=( a209a ) or ( a210a );
 a6507a <=( a211a ) or ( a6506a );
 a6508a <=( a6507a ) or ( a6502a );
 a6509a <=( a6508a ) or ( a6499a );
 a6512a <=( a207a ) or ( a208a );
 a6515a <=( a205a ) or ( a206a );
 a6516a <=( a6515a ) or ( a6512a );
 a6519a <=( a203a ) or ( a204a );
 a6523a <=( a200a ) or ( a201a );
 a6524a <=( a202a ) or ( a6523a );
 a6525a <=( a6524a ) or ( a6519a );
 a6526a <=( a6525a ) or ( a6516a );
 a6527a <=( a6526a ) or ( a6509a );
 a6530a <=( a198a ) or ( a199a );
 a6533a <=( a196a ) or ( a197a );
 a6534a <=( a6533a ) or ( a6530a );
 a6537a <=( a194a ) or ( a195a );
 a6541a <=( a191a ) or ( a192a );
 a6542a <=( a193a ) or ( a6541a );
 a6543a <=( a6542a ) or ( a6537a );
 a6544a <=( a6543a ) or ( a6534a );
 a6547a <=( a189a ) or ( a190a );
 a6550a <=( a187a ) or ( a188a );
 a6551a <=( a6550a ) or ( a6547a );
 a6554a <=( a185a ) or ( a186a );
 a6558a <=( a182a ) or ( a183a );
 a6559a <=( a184a ) or ( a6558a );
 a6560a <=( a6559a ) or ( a6554a );
 a6561a <=( a6560a ) or ( a6551a );
 a6562a <=( a6561a ) or ( a6544a );
 a6563a <=( a6562a ) or ( a6527a );
 a6566a <=( a180a ) or ( a181a );
 a6569a <=( a178a ) or ( a179a );
 a6570a <=( a6569a ) or ( a6566a );
 a6573a <=( a176a ) or ( a177a );
 a6577a <=( a173a ) or ( a174a );
 a6578a <=( a175a ) or ( a6577a );
 a6579a <=( a6578a ) or ( a6573a );
 a6580a <=( a6579a ) or ( a6570a );
 a6583a <=( a171a ) or ( a172a );
 a6586a <=( a169a ) or ( a170a );
 a6587a <=( a6586a ) or ( a6583a );
 a6590a <=( a167a ) or ( a168a );
 a6594a <=( a164a ) or ( a165a );
 a6595a <=( a166a ) or ( a6594a );
 a6596a <=( a6595a ) or ( a6590a );
 a6597a <=( a6596a ) or ( a6587a );
 a6598a <=( a6597a ) or ( a6580a );
 a6601a <=( a162a ) or ( a163a );
 a6604a <=( a160a ) or ( a161a );
 a6605a <=( a6604a ) or ( a6601a );
 a6608a <=( a158a ) or ( a159a );
 a6612a <=( a155a ) or ( a156a );
 a6613a <=( a157a ) or ( a6612a );
 a6614a <=( a6613a ) or ( a6608a );
 a6615a <=( a6614a ) or ( a6605a );
 a6618a <=( a153a ) or ( a154a );
 a6621a <=( a151a ) or ( a152a );
 a6622a <=( a6621a ) or ( a6618a );
 a6625a <=( a149a ) or ( a150a );
 a6629a <=( a146a ) or ( a147a );
 a6630a <=( a148a ) or ( a6629a );
 a6631a <=( a6630a ) or ( a6625a );
 a6632a <=( a6631a ) or ( a6622a );
 a6633a <=( a6632a ) or ( a6615a );
 a6634a <=( a6633a ) or ( a6598a );
 a6635a <=( a6634a ) or ( a6563a );
 a6636a <=( a6635a ) or ( a6492a );
 a6639a <=( a144a ) or ( a145a );
 a6642a <=( a142a ) or ( a143a );
 a6643a <=( a6642a ) or ( a6639a );
 a6646a <=( a140a ) or ( a141a );
 a6650a <=( a137a ) or ( a138a );
 a6651a <=( a139a ) or ( a6650a );
 a6652a <=( a6651a ) or ( a6646a );
 a6653a <=( a6652a ) or ( a6643a );
 a6656a <=( a135a ) or ( a136a );
 a6659a <=( a133a ) or ( a134a );
 a6660a <=( a6659a ) or ( a6656a );
 a6663a <=( a131a ) or ( a132a );
 a6667a <=( a128a ) or ( a129a );
 a6668a <=( a130a ) or ( a6667a );
 a6669a <=( a6668a ) or ( a6663a );
 a6670a <=( a6669a ) or ( a6660a );
 a6671a <=( a6670a ) or ( a6653a );
 a6674a <=( a126a ) or ( a127a );
 a6677a <=( a124a ) or ( a125a );
 a6678a <=( a6677a ) or ( a6674a );
 a6681a <=( a122a ) or ( a123a );
 a6685a <=( a119a ) or ( a120a );
 a6686a <=( a121a ) or ( a6685a );
 a6687a <=( a6686a ) or ( a6681a );
 a6688a <=( a6687a ) or ( a6678a );
 a6691a <=( a117a ) or ( a118a );
 a6694a <=( a115a ) or ( a116a );
 a6695a <=( a6694a ) or ( a6691a );
 a6698a <=( a113a ) or ( a114a );
 a6702a <=( a110a ) or ( a111a );
 a6703a <=( a112a ) or ( a6702a );
 a6704a <=( a6703a ) or ( a6698a );
 a6705a <=( a6704a ) or ( a6695a );
 a6706a <=( a6705a ) or ( a6688a );
 a6707a <=( a6706a ) or ( a6671a );
 a6710a <=( a108a ) or ( a109a );
 a6713a <=( a106a ) or ( a107a );
 a6714a <=( a6713a ) or ( a6710a );
 a6717a <=( a104a ) or ( a105a );
 a6721a <=( a101a ) or ( a102a );
 a6722a <=( a103a ) or ( a6721a );
 a6723a <=( a6722a ) or ( a6717a );
 a6724a <=( a6723a ) or ( a6714a );
 a6727a <=( a99a ) or ( a100a );
 a6730a <=( a97a ) or ( a98a );
 a6731a <=( a6730a ) or ( a6727a );
 a6734a <=( a95a ) or ( a96a );
 a6738a <=( a92a ) or ( a93a );
 a6739a <=( a94a ) or ( a6738a );
 a6740a <=( a6739a ) or ( a6734a );
 a6741a <=( a6740a ) or ( a6731a );
 a6742a <=( a6741a ) or ( a6724a );
 a6745a <=( a90a ) or ( a91a );
 a6748a <=( a88a ) or ( a89a );
 a6749a <=( a6748a ) or ( a6745a );
 a6752a <=( a86a ) or ( a87a );
 a6756a <=( a83a ) or ( a84a );
 a6757a <=( a85a ) or ( a6756a );
 a6758a <=( a6757a ) or ( a6752a );
 a6759a <=( a6758a ) or ( a6749a );
 a6762a <=( a81a ) or ( a82a );
 a6765a <=( a79a ) or ( a80a );
 a6766a <=( a6765a ) or ( a6762a );
 a6769a <=( a77a ) or ( a78a );
 a6773a <=( a74a ) or ( a75a );
 a6774a <=( a76a ) or ( a6773a );
 a6775a <=( a6774a ) or ( a6769a );
 a6776a <=( a6775a ) or ( a6766a );
 a6777a <=( a6776a ) or ( a6759a );
 a6778a <=( a6777a ) or ( a6742a );
 a6779a <=( a6778a ) or ( a6707a );
 a6782a <=( a72a ) or ( a73a );
 a6785a <=( a70a ) or ( a71a );
 a6786a <=( a6785a ) or ( a6782a );
 a6789a <=( a68a ) or ( a69a );
 a6793a <=( a65a ) or ( a66a );
 a6794a <=( a67a ) or ( a6793a );
 a6795a <=( a6794a ) or ( a6789a );
 a6796a <=( a6795a ) or ( a6786a );
 a6799a <=( a63a ) or ( a64a );
 a6802a <=( a61a ) or ( a62a );
 a6803a <=( a6802a ) or ( a6799a );
 a6806a <=( a59a ) or ( a60a );
 a6810a <=( a56a ) or ( a57a );
 a6811a <=( a58a ) or ( a6810a );
 a6812a <=( a6811a ) or ( a6806a );
 a6813a <=( a6812a ) or ( a6803a );
 a6814a <=( a6813a ) or ( a6796a );
 a6817a <=( a54a ) or ( a55a );
 a6820a <=( a52a ) or ( a53a );
 a6821a <=( a6820a ) or ( a6817a );
 a6824a <=( a50a ) or ( a51a );
 a6828a <=( a47a ) or ( a48a );
 a6829a <=( a49a ) or ( a6828a );
 a6830a <=( a6829a ) or ( a6824a );
 a6831a <=( a6830a ) or ( a6821a );
 a6834a <=( a45a ) or ( a46a );
 a6837a <=( a43a ) or ( a44a );
 a6838a <=( a6837a ) or ( a6834a );
 a6841a <=( a41a ) or ( a42a );
 a6845a <=( a38a ) or ( a39a );
 a6846a <=( a40a ) or ( a6845a );
 a6847a <=( a6846a ) or ( a6841a );
 a6848a <=( a6847a ) or ( a6838a );
 a6849a <=( a6848a ) or ( a6831a );
 a6850a <=( a6849a ) or ( a6814a );
 a6853a <=( a36a ) or ( a37a );
 a6856a <=( a34a ) or ( a35a );
 a6857a <=( a6856a ) or ( a6853a );
 a6860a <=( a32a ) or ( a33a );
 a6864a <=( a29a ) or ( a30a );
 a6865a <=( a31a ) or ( a6864a );
 a6866a <=( a6865a ) or ( a6860a );
 a6867a <=( a6866a ) or ( a6857a );
 a6870a <=( a27a ) or ( a28a );
 a6873a <=( a25a ) or ( a26a );
 a6874a <=( a6873a ) or ( a6870a );
 a6877a <=( a23a ) or ( a24a );
 a6881a <=( a20a ) or ( a21a );
 a6882a <=( a22a ) or ( a6881a );
 a6883a <=( a6882a ) or ( a6877a );
 a6884a <=( a6883a ) or ( a6874a );
 a6885a <=( a6884a ) or ( a6867a );
 a6888a <=( a18a ) or ( a19a );
 a6891a <=( a16a ) or ( a17a );
 a6892a <=( a6891a ) or ( a6888a );
 a6895a <=( a14a ) or ( a15a );
 a6899a <=( a11a ) or ( a12a );
 a6900a <=( a13a ) or ( a6899a );
 a6901a <=( a6900a ) or ( a6895a );
 a6902a <=( a6901a ) or ( a6892a );
 a6905a <=( a9a ) or ( a10a );
 a6909a <=( a6a ) or ( a7a );
 a6910a <=( a8a ) or ( a6909a );
 a6911a <=( a6910a ) or ( a6905a );
 a6914a <=( a4a ) or ( a5a );
 a6918a <=( a1a ) or ( a2a );
 a6919a <=( a3a ) or ( a6918a );
 a6920a <=( a6919a ) or ( a6914a );
 a6921a <=( a6920a ) or ( a6911a );
 a6922a <=( a6921a ) or ( a6902a );
 a6923a <=( a6922a ) or ( a6885a );
 a6924a <=( a6923a ) or ( a6850a );
 a6925a <=( a6924a ) or ( a6779a );
 a6926a <=( a6925a ) or ( a6636a );
 a6927a <=( a6926a ) or ( a6349a );
 a6928a <=( a6927a ) or ( a5772a );
 a6932a <=( (not A202)  and  (not A201) );
 a6933a <=( A169  and  a6932a );
 a6937a <=( A301  and  A235 );
 a6938a <=( (not A203)  and  a6937a );
 a6942a <=( (not A202)  and  (not A201) );
 a6943a <=( A169  and  a6942a );
 a6947a <=( A268  and  A235 );
 a6948a <=( (not A203)  and  a6947a );
 a6952a <=( (not A200)  and  (not A199) );
 a6953a <=( A169  and  a6952a );
 a6957a <=( A301  and  A235 );
 a6958a <=( (not A202)  and  a6957a );
 a6962a <=( (not A200)  and  (not A199) );
 a6963a <=( A169  and  a6962a );
 a6967a <=( A268  and  A235 );
 a6968a <=( (not A202)  and  a6967a );
 a6972a <=( (not A166)  and  (not A167) );
 a6973a <=( (not A169)  and  a6972a );
 a6977a <=( A301  and  A235 );
 a6978a <=( A202  and  a6977a );
 a6982a <=( (not A166)  and  (not A167) );
 a6983a <=( (not A169)  and  a6982a );
 a6987a <=( A268  and  A235 );
 a6988a <=( A202  and  a6987a );
 a6992a <=( (not A168)  and  (not A169) );
 a6993a <=( (not A170)  and  a6992a );
 a6997a <=( A301  and  A235 );
 a6998a <=( A202  and  a6997a );
 a7002a <=( (not A168)  and  (not A169) );
 a7003a <=( (not A170)  and  a7002a );
 a7007a <=( A268  and  A235 );
 a7008a <=( A202  and  a7007a );
 a7012a <=( (not A201)  and  A166 );
 a7013a <=( A168  and  a7012a );
 a7016a <=( (not A203)  and  (not A202) );
 a7019a <=( A301  and  A235 );
 a7020a <=( a7019a  and  a7016a );
 a7024a <=( (not A201)  and  A166 );
 a7025a <=( A168  and  a7024a );
 a7028a <=( (not A203)  and  (not A202) );
 a7031a <=( A268  and  A235 );
 a7032a <=( a7031a  and  a7028a );
 a7036a <=( (not A199)  and  A166 );
 a7037a <=( A168  and  a7036a );
 a7040a <=( (not A202)  and  (not A200) );
 a7043a <=( A301  and  A235 );
 a7044a <=( a7043a  and  a7040a );
 a7048a <=( (not A199)  and  A166 );
 a7049a <=( A168  and  a7048a );
 a7052a <=( (not A202)  and  (not A200) );
 a7055a <=( A268  and  A235 );
 a7056a <=( a7055a  and  a7052a );
 a7060a <=( (not A201)  and  A167 );
 a7061a <=( A168  and  a7060a );
 a7064a <=( (not A203)  and  (not A202) );
 a7067a <=( A301  and  A235 );
 a7068a <=( a7067a  and  a7064a );
 a7072a <=( (not A201)  and  A167 );
 a7073a <=( A168  and  a7072a );
 a7076a <=( (not A203)  and  (not A202) );
 a7079a <=( A268  and  A235 );
 a7080a <=( a7079a  and  a7076a );
 a7084a <=( (not A199)  and  A167 );
 a7085a <=( A168  and  a7084a );
 a7088a <=( (not A202)  and  (not A200) );
 a7091a <=( A301  and  A235 );
 a7092a <=( a7091a  and  a7088a );
 a7096a <=( (not A199)  and  A167 );
 a7097a <=( A168  and  a7096a );
 a7100a <=( (not A202)  and  (not A200) );
 a7103a <=( A268  and  A235 );
 a7104a <=( a7103a  and  a7100a );
 a7108a <=( (not A202)  and  (not A201) );
 a7109a <=( A169  and  a7108a );
 a7112a <=( A235  and  (not A203) );
 a7115a <=( A300  and  A299 );
 a7116a <=( a7115a  and  a7112a );
 a7120a <=( (not A202)  and  (not A201) );
 a7121a <=( A169  and  a7120a );
 a7124a <=( A235  and  (not A203) );
 a7127a <=( A300  and  A298 );
 a7128a <=( a7127a  and  a7124a );
 a7132a <=( (not A202)  and  (not A201) );
 a7133a <=( A169  and  a7132a );
 a7136a <=( A235  and  (not A203) );
 a7139a <=( A267  and  A265 );
 a7140a <=( a7139a  and  a7136a );
 a7144a <=( (not A202)  and  (not A201) );
 a7145a <=( A169  and  a7144a );
 a7148a <=( A235  and  (not A203) );
 a7151a <=( A267  and  A266 );
 a7152a <=( a7151a  and  a7148a );
 a7156a <=( (not A202)  and  (not A201) );
 a7157a <=( A169  and  a7156a );
 a7160a <=( A232  and  (not A203) );
 a7163a <=( A301  and  A234 );
 a7164a <=( a7163a  and  a7160a );
 a7168a <=( (not A202)  and  (not A201) );
 a7169a <=( A169  and  a7168a );
 a7172a <=( A232  and  (not A203) );
 a7175a <=( A268  and  A234 );
 a7176a <=( a7175a  and  a7172a );
 a7180a <=( (not A202)  and  (not A201) );
 a7181a <=( A169  and  a7180a );
 a7184a <=( A233  and  (not A203) );
 a7187a <=( A301  and  A234 );
 a7188a <=( a7187a  and  a7184a );
 a7192a <=( (not A202)  and  (not A201) );
 a7193a <=( A169  and  a7192a );
 a7196a <=( A233  and  (not A203) );
 a7199a <=( A268  and  A234 );
 a7200a <=( a7199a  and  a7196a );
 a7204a <=( A200  and  A199 );
 a7205a <=( A169  and  a7204a );
 a7208a <=( (not A202)  and  (not A201) );
 a7211a <=( A301  and  A235 );
 a7212a <=( a7211a  and  a7208a );
 a7216a <=( A200  and  A199 );
 a7217a <=( A169  and  a7216a );
 a7220a <=( (not A202)  and  (not A201) );
 a7223a <=( A268  and  A235 );
 a7224a <=( a7223a  and  a7220a );
 a7228a <=( (not A200)  and  (not A199) );
 a7229a <=( A169  and  a7228a );
 a7232a <=( A235  and  (not A202) );
 a7235a <=( A300  and  A299 );
 a7236a <=( a7235a  and  a7232a );
 a7240a <=( (not A200)  and  (not A199) );
 a7241a <=( A169  and  a7240a );
 a7244a <=( A235  and  (not A202) );
 a7247a <=( A300  and  A298 );
 a7248a <=( a7247a  and  a7244a );
 a7252a <=( (not A200)  and  (not A199) );
 a7253a <=( A169  and  a7252a );
 a7256a <=( A235  and  (not A202) );
 a7259a <=( A267  and  A265 );
 a7260a <=( a7259a  and  a7256a );
 a7264a <=( (not A200)  and  (not A199) );
 a7265a <=( A169  and  a7264a );
 a7268a <=( A235  and  (not A202) );
 a7271a <=( A267  and  A266 );
 a7272a <=( a7271a  and  a7268a );
 a7276a <=( (not A200)  and  (not A199) );
 a7277a <=( A169  and  a7276a );
 a7280a <=( A232  and  (not A202) );
 a7283a <=( A301  and  A234 );
 a7284a <=( a7283a  and  a7280a );
 a7288a <=( (not A200)  and  (not A199) );
 a7289a <=( A169  and  a7288a );
 a7292a <=( A232  and  (not A202) );
 a7295a <=( A268  and  A234 );
 a7296a <=( a7295a  and  a7292a );
 a7300a <=( (not A200)  and  (not A199) );
 a7301a <=( A169  and  a7300a );
 a7304a <=( A233  and  (not A202) );
 a7307a <=( A301  and  A234 );
 a7308a <=( a7307a  and  a7304a );
 a7312a <=( (not A200)  and  (not A199) );
 a7313a <=( A169  and  a7312a );
 a7316a <=( A233  and  (not A202) );
 a7319a <=( A268  and  A234 );
 a7320a <=( a7319a  and  a7316a );
 a7324a <=( (not A166)  and  (not A167) );
 a7325a <=( (not A169)  and  a7324a );
 a7328a <=( A235  and  A202 );
 a7331a <=( A300  and  A299 );
 a7332a <=( a7331a  and  a7328a );
 a7336a <=( (not A166)  and  (not A167) );
 a7337a <=( (not A169)  and  a7336a );
 a7340a <=( A235  and  A202 );
 a7343a <=( A300  and  A298 );
 a7344a <=( a7343a  and  a7340a );
 a7348a <=( (not A166)  and  (not A167) );
 a7349a <=( (not A169)  and  a7348a );
 a7352a <=( A235  and  A202 );
 a7355a <=( A267  and  A265 );
 a7356a <=( a7355a  and  a7352a );
 a7360a <=( (not A166)  and  (not A167) );
 a7361a <=( (not A169)  and  a7360a );
 a7364a <=( A235  and  A202 );
 a7367a <=( A267  and  A266 );
 a7368a <=( a7367a  and  a7364a );
 a7372a <=( (not A166)  and  (not A167) );
 a7373a <=( (not A169)  and  a7372a );
 a7376a <=( A232  and  A202 );
 a7379a <=( A301  and  A234 );
 a7380a <=( a7379a  and  a7376a );
 a7384a <=( (not A166)  and  (not A167) );
 a7385a <=( (not A169)  and  a7384a );
 a7388a <=( A232  and  A202 );
 a7391a <=( A268  and  A234 );
 a7392a <=( a7391a  and  a7388a );
 a7396a <=( (not A166)  and  (not A167) );
 a7397a <=( (not A169)  and  a7396a );
 a7400a <=( A233  and  A202 );
 a7403a <=( A301  and  A234 );
 a7404a <=( a7403a  and  a7400a );
 a7408a <=( (not A166)  and  (not A167) );
 a7409a <=( (not A169)  and  a7408a );
 a7412a <=( A233  and  A202 );
 a7415a <=( A268  and  A234 );
 a7416a <=( a7415a  and  a7412a );
 a7420a <=( (not A166)  and  (not A167) );
 a7421a <=( (not A169)  and  a7420a );
 a7424a <=( A201  and  A199 );
 a7427a <=( A301  and  A235 );
 a7428a <=( a7427a  and  a7424a );
 a7432a <=( (not A166)  and  (not A167) );
 a7433a <=( (not A169)  and  a7432a );
 a7436a <=( A201  and  A199 );
 a7439a <=( A268  and  A235 );
 a7440a <=( a7439a  and  a7436a );
 a7444a <=( (not A166)  and  (not A167) );
 a7445a <=( (not A169)  and  a7444a );
 a7448a <=( A201  and  A200 );
 a7451a <=( A301  and  A235 );
 a7452a <=( a7451a  and  a7448a );
 a7456a <=( (not A166)  and  (not A167) );
 a7457a <=( (not A169)  and  a7456a );
 a7460a <=( A201  and  A200 );
 a7463a <=( A268  and  A235 );
 a7464a <=( a7463a  and  a7460a );
 a7468a <=( A167  and  (not A168) );
 a7469a <=( (not A169)  and  a7468a );
 a7472a <=( A202  and  A166 );
 a7475a <=( A301  and  A235 );
 a7476a <=( a7475a  and  a7472a );
 a7480a <=( A167  and  (not A168) );
 a7481a <=( (not A169)  and  a7480a );
 a7484a <=( A202  and  A166 );
 a7487a <=( A268  and  A235 );
 a7488a <=( a7487a  and  a7484a );
 a7492a <=( (not A168)  and  (not A169) );
 a7493a <=( (not A170)  and  a7492a );
 a7496a <=( A235  and  A202 );
 a7499a <=( A300  and  A299 );
 a7500a <=( a7499a  and  a7496a );
 a7504a <=( (not A168)  and  (not A169) );
 a7505a <=( (not A170)  and  a7504a );
 a7508a <=( A235  and  A202 );
 a7511a <=( A300  and  A298 );
 a7512a <=( a7511a  and  a7508a );
 a7516a <=( (not A168)  and  (not A169) );
 a7517a <=( (not A170)  and  a7516a );
 a7520a <=( A235  and  A202 );
 a7523a <=( A267  and  A265 );
 a7524a <=( a7523a  and  a7520a );
 a7528a <=( (not A168)  and  (not A169) );
 a7529a <=( (not A170)  and  a7528a );
 a7532a <=( A235  and  A202 );
 a7535a <=( A267  and  A266 );
 a7536a <=( a7535a  and  a7532a );
 a7540a <=( (not A168)  and  (not A169) );
 a7541a <=( (not A170)  and  a7540a );
 a7544a <=( A232  and  A202 );
 a7547a <=( A301  and  A234 );
 a7548a <=( a7547a  and  a7544a );
 a7552a <=( (not A168)  and  (not A169) );
 a7553a <=( (not A170)  and  a7552a );
 a7556a <=( A232  and  A202 );
 a7559a <=( A268  and  A234 );
 a7560a <=( a7559a  and  a7556a );
 a7564a <=( (not A168)  and  (not A169) );
 a7565a <=( (not A170)  and  a7564a );
 a7568a <=( A233  and  A202 );
 a7571a <=( A301  and  A234 );
 a7572a <=( a7571a  and  a7568a );
 a7576a <=( (not A168)  and  (not A169) );
 a7577a <=( (not A170)  and  a7576a );
 a7580a <=( A233  and  A202 );
 a7583a <=( A268  and  A234 );
 a7584a <=( a7583a  and  a7580a );
 a7588a <=( (not A168)  and  (not A169) );
 a7589a <=( (not A170)  and  a7588a );
 a7592a <=( A201  and  A199 );
 a7595a <=( A301  and  A235 );
 a7596a <=( a7595a  and  a7592a );
 a7600a <=( (not A168)  and  (not A169) );
 a7601a <=( (not A170)  and  a7600a );
 a7604a <=( A201  and  A199 );
 a7607a <=( A268  and  A235 );
 a7608a <=( a7607a  and  a7604a );
 a7612a <=( (not A168)  and  (not A169) );
 a7613a <=( (not A170)  and  a7612a );
 a7616a <=( A201  and  A200 );
 a7619a <=( A301  and  A235 );
 a7620a <=( a7619a  and  a7616a );
 a7624a <=( (not A168)  and  (not A169) );
 a7625a <=( (not A170)  and  a7624a );
 a7628a <=( A201  and  A200 );
 a7631a <=( A268  and  A235 );
 a7632a <=( a7631a  and  a7628a );
 a7635a <=( A166  and  A168 );
 a7638a <=( (not A202)  and  (not A201) );
 a7639a <=( a7638a  and  a7635a );
 a7642a <=( A235  and  (not A203) );
 a7645a <=( A300  and  A299 );
 a7646a <=( a7645a  and  a7642a );
 a7649a <=( A166  and  A168 );
 a7652a <=( (not A202)  and  (not A201) );
 a7653a <=( a7652a  and  a7649a );
 a7656a <=( A235  and  (not A203) );
 a7659a <=( A300  and  A298 );
 a7660a <=( a7659a  and  a7656a );
 a7663a <=( A166  and  A168 );
 a7666a <=( (not A202)  and  (not A201) );
 a7667a <=( a7666a  and  a7663a );
 a7670a <=( A235  and  (not A203) );
 a7673a <=( A267  and  A265 );
 a7674a <=( a7673a  and  a7670a );
 a7677a <=( A166  and  A168 );
 a7680a <=( (not A202)  and  (not A201) );
 a7681a <=( a7680a  and  a7677a );
 a7684a <=( A235  and  (not A203) );
 a7687a <=( A267  and  A266 );
 a7688a <=( a7687a  and  a7684a );
 a7691a <=( A166  and  A168 );
 a7694a <=( (not A202)  and  (not A201) );
 a7695a <=( a7694a  and  a7691a );
 a7698a <=( A232  and  (not A203) );
 a7701a <=( A301  and  A234 );
 a7702a <=( a7701a  and  a7698a );
 a7705a <=( A166  and  A168 );
 a7708a <=( (not A202)  and  (not A201) );
 a7709a <=( a7708a  and  a7705a );
 a7712a <=( A232  and  (not A203) );
 a7715a <=( A268  and  A234 );
 a7716a <=( a7715a  and  a7712a );
 a7719a <=( A166  and  A168 );
 a7722a <=( (not A202)  and  (not A201) );
 a7723a <=( a7722a  and  a7719a );
 a7726a <=( A233  and  (not A203) );
 a7729a <=( A301  and  A234 );
 a7730a <=( a7729a  and  a7726a );
 a7733a <=( A166  and  A168 );
 a7736a <=( (not A202)  and  (not A201) );
 a7737a <=( a7736a  and  a7733a );
 a7740a <=( A233  and  (not A203) );
 a7743a <=( A268  and  A234 );
 a7744a <=( a7743a  and  a7740a );
 a7747a <=( A166  and  A168 );
 a7750a <=( A200  and  A199 );
 a7751a <=( a7750a  and  a7747a );
 a7754a <=( (not A202)  and  (not A201) );
 a7757a <=( A301  and  A235 );
 a7758a <=( a7757a  and  a7754a );
 a7761a <=( A166  and  A168 );
 a7764a <=( A200  and  A199 );
 a7765a <=( a7764a  and  a7761a );
 a7768a <=( (not A202)  and  (not A201) );
 a7771a <=( A268  and  A235 );
 a7772a <=( a7771a  and  a7768a );
 a7775a <=( A166  and  A168 );
 a7778a <=( (not A200)  and  (not A199) );
 a7779a <=( a7778a  and  a7775a );
 a7782a <=( A235  and  (not A202) );
 a7785a <=( A300  and  A299 );
 a7786a <=( a7785a  and  a7782a );
 a7789a <=( A166  and  A168 );
 a7792a <=( (not A200)  and  (not A199) );
 a7793a <=( a7792a  and  a7789a );
 a7796a <=( A235  and  (not A202) );
 a7799a <=( A300  and  A298 );
 a7800a <=( a7799a  and  a7796a );
 a7803a <=( A166  and  A168 );
 a7806a <=( (not A200)  and  (not A199) );
 a7807a <=( a7806a  and  a7803a );
 a7810a <=( A235  and  (not A202) );
 a7813a <=( A267  and  A265 );
 a7814a <=( a7813a  and  a7810a );
 a7817a <=( A166  and  A168 );
 a7820a <=( (not A200)  and  (not A199) );
 a7821a <=( a7820a  and  a7817a );
 a7824a <=( A235  and  (not A202) );
 a7827a <=( A267  and  A266 );
 a7828a <=( a7827a  and  a7824a );
 a7831a <=( A166  and  A168 );
 a7834a <=( (not A200)  and  (not A199) );
 a7835a <=( a7834a  and  a7831a );
 a7838a <=( A232  and  (not A202) );
 a7841a <=( A301  and  A234 );
 a7842a <=( a7841a  and  a7838a );
 a7845a <=( A166  and  A168 );
 a7848a <=( (not A200)  and  (not A199) );
 a7849a <=( a7848a  and  a7845a );
 a7852a <=( A232  and  (not A202) );
 a7855a <=( A268  and  A234 );
 a7856a <=( a7855a  and  a7852a );
 a7859a <=( A166  and  A168 );
 a7862a <=( (not A200)  and  (not A199) );
 a7863a <=( a7862a  and  a7859a );
 a7866a <=( A233  and  (not A202) );
 a7869a <=( A301  and  A234 );
 a7870a <=( a7869a  and  a7866a );
 a7873a <=( A166  and  A168 );
 a7876a <=( (not A200)  and  (not A199) );
 a7877a <=( a7876a  and  a7873a );
 a7880a <=( A233  and  (not A202) );
 a7883a <=( A268  and  A234 );
 a7884a <=( a7883a  and  a7880a );
 a7887a <=( A167  and  A168 );
 a7890a <=( (not A202)  and  (not A201) );
 a7891a <=( a7890a  and  a7887a );
 a7894a <=( A235  and  (not A203) );
 a7897a <=( A300  and  A299 );
 a7898a <=( a7897a  and  a7894a );
 a7901a <=( A167  and  A168 );
 a7904a <=( (not A202)  and  (not A201) );
 a7905a <=( a7904a  and  a7901a );
 a7908a <=( A235  and  (not A203) );
 a7911a <=( A300  and  A298 );
 a7912a <=( a7911a  and  a7908a );
 a7915a <=( A167  and  A168 );
 a7918a <=( (not A202)  and  (not A201) );
 a7919a <=( a7918a  and  a7915a );
 a7922a <=( A235  and  (not A203) );
 a7925a <=( A267  and  A265 );
 a7926a <=( a7925a  and  a7922a );
 a7929a <=( A167  and  A168 );
 a7932a <=( (not A202)  and  (not A201) );
 a7933a <=( a7932a  and  a7929a );
 a7936a <=( A235  and  (not A203) );
 a7939a <=( A267  and  A266 );
 a7940a <=( a7939a  and  a7936a );
 a7943a <=( A167  and  A168 );
 a7946a <=( (not A202)  and  (not A201) );
 a7947a <=( a7946a  and  a7943a );
 a7950a <=( A232  and  (not A203) );
 a7953a <=( A301  and  A234 );
 a7954a <=( a7953a  and  a7950a );
 a7957a <=( A167  and  A168 );
 a7960a <=( (not A202)  and  (not A201) );
 a7961a <=( a7960a  and  a7957a );
 a7964a <=( A232  and  (not A203) );
 a7967a <=( A268  and  A234 );
 a7968a <=( a7967a  and  a7964a );
 a7971a <=( A167  and  A168 );
 a7974a <=( (not A202)  and  (not A201) );
 a7975a <=( a7974a  and  a7971a );
 a7978a <=( A233  and  (not A203) );
 a7981a <=( A301  and  A234 );
 a7982a <=( a7981a  and  a7978a );
 a7985a <=( A167  and  A168 );
 a7988a <=( (not A202)  and  (not A201) );
 a7989a <=( a7988a  and  a7985a );
 a7992a <=( A233  and  (not A203) );
 a7995a <=( A268  and  A234 );
 a7996a <=( a7995a  and  a7992a );
 a7999a <=( A167  and  A168 );
 a8002a <=( A200  and  A199 );
 a8003a <=( a8002a  and  a7999a );
 a8006a <=( (not A202)  and  (not A201) );
 a8009a <=( A301  and  A235 );
 a8010a <=( a8009a  and  a8006a );
 a8013a <=( A167  and  A168 );
 a8016a <=( A200  and  A199 );
 a8017a <=( a8016a  and  a8013a );
 a8020a <=( (not A202)  and  (not A201) );
 a8023a <=( A268  and  A235 );
 a8024a <=( a8023a  and  a8020a );
 a8027a <=( A167  and  A168 );
 a8030a <=( (not A200)  and  (not A199) );
 a8031a <=( a8030a  and  a8027a );
 a8034a <=( A235  and  (not A202) );
 a8037a <=( A300  and  A299 );
 a8038a <=( a8037a  and  a8034a );
 a8041a <=( A167  and  A168 );
 a8044a <=( (not A200)  and  (not A199) );
 a8045a <=( a8044a  and  a8041a );
 a8048a <=( A235  and  (not A202) );
 a8051a <=( A300  and  A298 );
 a8052a <=( a8051a  and  a8048a );
 a8055a <=( A167  and  A168 );
 a8058a <=( (not A200)  and  (not A199) );
 a8059a <=( a8058a  and  a8055a );
 a8062a <=( A235  and  (not A202) );
 a8065a <=( A267  and  A265 );
 a8066a <=( a8065a  and  a8062a );
 a8069a <=( A167  and  A168 );
 a8072a <=( (not A200)  and  (not A199) );
 a8073a <=( a8072a  and  a8069a );
 a8076a <=( A235  and  (not A202) );
 a8079a <=( A267  and  A266 );
 a8080a <=( a8079a  and  a8076a );
 a8083a <=( A167  and  A168 );
 a8086a <=( (not A200)  and  (not A199) );
 a8087a <=( a8086a  and  a8083a );
 a8090a <=( A232  and  (not A202) );
 a8093a <=( A301  and  A234 );
 a8094a <=( a8093a  and  a8090a );
 a8097a <=( A167  and  A168 );
 a8100a <=( (not A200)  and  (not A199) );
 a8101a <=( a8100a  and  a8097a );
 a8104a <=( A232  and  (not A202) );
 a8107a <=( A268  and  A234 );
 a8108a <=( a8107a  and  a8104a );
 a8111a <=( A167  and  A168 );
 a8114a <=( (not A200)  and  (not A199) );
 a8115a <=( a8114a  and  a8111a );
 a8118a <=( A233  and  (not A202) );
 a8121a <=( A301  and  A234 );
 a8122a <=( a8121a  and  a8118a );
 a8125a <=( A167  and  A168 );
 a8128a <=( (not A200)  and  (not A199) );
 a8129a <=( a8128a  and  a8125a );
 a8132a <=( A233  and  (not A202) );
 a8135a <=( A268  and  A234 );
 a8136a <=( a8135a  and  a8132a );
 a8139a <=( A167  and  A170 );
 a8142a <=( (not A201)  and  (not A166) );
 a8143a <=( a8142a  and  a8139a );
 a8146a <=( (not A203)  and  (not A202) );
 a8149a <=( A301  and  A235 );
 a8150a <=( a8149a  and  a8146a );
 a8153a <=( A167  and  A170 );
 a8156a <=( (not A201)  and  (not A166) );
 a8157a <=( a8156a  and  a8153a );
 a8160a <=( (not A203)  and  (not A202) );
 a8163a <=( A268  and  A235 );
 a8164a <=( a8163a  and  a8160a );
 a8167a <=( A167  and  A170 );
 a8170a <=( (not A199)  and  (not A166) );
 a8171a <=( a8170a  and  a8167a );
 a8174a <=( (not A202)  and  (not A200) );
 a8177a <=( A301  and  A235 );
 a8178a <=( a8177a  and  a8174a );
 a8181a <=( A167  and  A170 );
 a8184a <=( (not A199)  and  (not A166) );
 a8185a <=( a8184a  and  a8181a );
 a8188a <=( (not A202)  and  (not A200) );
 a8191a <=( A268  and  A235 );
 a8192a <=( a8191a  and  a8188a );
 a8195a <=( (not A167)  and  A170 );
 a8198a <=( (not A201)  and  A166 );
 a8199a <=( a8198a  and  a8195a );
 a8202a <=( (not A203)  and  (not A202) );
 a8205a <=( A301  and  A235 );
 a8206a <=( a8205a  and  a8202a );
 a8209a <=( (not A167)  and  A170 );
 a8212a <=( (not A201)  and  A166 );
 a8213a <=( a8212a  and  a8209a );
 a8216a <=( (not A203)  and  (not A202) );
 a8219a <=( A268  and  A235 );
 a8220a <=( a8219a  and  a8216a );
 a8223a <=( (not A167)  and  A170 );
 a8226a <=( (not A199)  and  A166 );
 a8227a <=( a8226a  and  a8223a );
 a8230a <=( (not A202)  and  (not A200) );
 a8233a <=( A301  and  A235 );
 a8234a <=( a8233a  and  a8230a );
 a8237a <=( (not A167)  and  A170 );
 a8240a <=( (not A199)  and  A166 );
 a8241a <=( a8240a  and  a8237a );
 a8244a <=( (not A202)  and  (not A200) );
 a8247a <=( A268  and  A235 );
 a8248a <=( a8247a  and  a8244a );
 a8251a <=( (not A201)  and  A169 );
 a8254a <=( (not A203)  and  (not A202) );
 a8255a <=( a8254a  and  a8251a );
 a8258a <=( A298  and  A235 );
 a8261a <=( A302  and  (not A299) );
 a8262a <=( a8261a  and  a8258a );
 a8265a <=( (not A201)  and  A169 );
 a8268a <=( (not A203)  and  (not A202) );
 a8269a <=( a8268a  and  a8265a );
 a8272a <=( (not A298)  and  A235 );
 a8275a <=( A302  and  A299 );
 a8276a <=( a8275a  and  a8272a );
 a8279a <=( (not A201)  and  A169 );
 a8282a <=( (not A203)  and  (not A202) );
 a8283a <=( a8282a  and  a8279a );
 a8286a <=( (not A265)  and  A235 );
 a8289a <=( A269  and  A266 );
 a8290a <=( a8289a  and  a8286a );
 a8293a <=( (not A201)  and  A169 );
 a8296a <=( (not A203)  and  (not A202) );
 a8297a <=( a8296a  and  a8293a );
 a8300a <=( A265  and  A235 );
 a8303a <=( A269  and  (not A266) );
 a8304a <=( a8303a  and  a8300a );
 a8307a <=( (not A201)  and  A169 );
 a8310a <=( (not A203)  and  (not A202) );
 a8311a <=( a8310a  and  a8307a );
 a8314a <=( A234  and  A232 );
 a8317a <=( A300  and  A299 );
 a8318a <=( a8317a  and  a8314a );
 a8321a <=( (not A201)  and  A169 );
 a8324a <=( (not A203)  and  (not A202) );
 a8325a <=( a8324a  and  a8321a );
 a8328a <=( A234  and  A232 );
 a8331a <=( A300  and  A298 );
 a8332a <=( a8331a  and  a8328a );
 a8335a <=( (not A201)  and  A169 );
 a8338a <=( (not A203)  and  (not A202) );
 a8339a <=( a8338a  and  a8335a );
 a8342a <=( A234  and  A232 );
 a8345a <=( A267  and  A265 );
 a8346a <=( a8345a  and  a8342a );
 a8349a <=( (not A201)  and  A169 );
 a8352a <=( (not A203)  and  (not A202) );
 a8353a <=( a8352a  and  a8349a );
 a8356a <=( A234  and  A232 );
 a8359a <=( A267  and  A266 );
 a8360a <=( a8359a  and  a8356a );
 a8363a <=( (not A201)  and  A169 );
 a8366a <=( (not A203)  and  (not A202) );
 a8367a <=( a8366a  and  a8363a );
 a8370a <=( A234  and  A233 );
 a8373a <=( A300  and  A299 );
 a8374a <=( a8373a  and  a8370a );
 a8377a <=( (not A201)  and  A169 );
 a8380a <=( (not A203)  and  (not A202) );
 a8381a <=( a8380a  and  a8377a );
 a8384a <=( A234  and  A233 );
 a8387a <=( A300  and  A298 );
 a8388a <=( a8387a  and  a8384a );
 a8391a <=( (not A201)  and  A169 );
 a8394a <=( (not A203)  and  (not A202) );
 a8395a <=( a8394a  and  a8391a );
 a8398a <=( A234  and  A233 );
 a8401a <=( A267  and  A265 );
 a8402a <=( a8401a  and  a8398a );
 a8405a <=( (not A201)  and  A169 );
 a8408a <=( (not A203)  and  (not A202) );
 a8409a <=( a8408a  and  a8405a );
 a8412a <=( A234  and  A233 );
 a8415a <=( A267  and  A266 );
 a8416a <=( a8415a  and  a8412a );
 a8419a <=( (not A201)  and  A169 );
 a8422a <=( (not A203)  and  (not A202) );
 a8423a <=( a8422a  and  a8419a );
 a8426a <=( A233  and  (not A232) );
 a8429a <=( A301  and  A236 );
 a8430a <=( a8429a  and  a8426a );
 a8433a <=( (not A201)  and  A169 );
 a8436a <=( (not A203)  and  (not A202) );
 a8437a <=( a8436a  and  a8433a );
 a8440a <=( A233  and  (not A232) );
 a8443a <=( A268  and  A236 );
 a8444a <=( a8443a  and  a8440a );
 a8447a <=( (not A201)  and  A169 );
 a8450a <=( (not A203)  and  (not A202) );
 a8451a <=( a8450a  and  a8447a );
 a8454a <=( (not A233)  and  A232 );
 a8457a <=( A301  and  A236 );
 a8458a <=( a8457a  and  a8454a );
 a8461a <=( (not A201)  and  A169 );
 a8464a <=( (not A203)  and  (not A202) );
 a8465a <=( a8464a  and  a8461a );
 a8468a <=( (not A233)  and  A232 );
 a8471a <=( A268  and  A236 );
 a8472a <=( a8471a  and  a8468a );
 a8475a <=( A199  and  A169 );
 a8478a <=( (not A201)  and  A200 );
 a8479a <=( a8478a  and  a8475a );
 a8482a <=( A235  and  (not A202) );
 a8485a <=( A300  and  A299 );
 a8486a <=( a8485a  and  a8482a );
 a8489a <=( A199  and  A169 );
 a8492a <=( (not A201)  and  A200 );
 a8493a <=( a8492a  and  a8489a );
 a8496a <=( A235  and  (not A202) );
 a8499a <=( A300  and  A298 );
 a8500a <=( a8499a  and  a8496a );
 a8503a <=( A199  and  A169 );
 a8506a <=( (not A201)  and  A200 );
 a8507a <=( a8506a  and  a8503a );
 a8510a <=( A235  and  (not A202) );
 a8513a <=( A267  and  A265 );
 a8514a <=( a8513a  and  a8510a );
 a8517a <=( A199  and  A169 );
 a8520a <=( (not A201)  and  A200 );
 a8521a <=( a8520a  and  a8517a );
 a8524a <=( A235  and  (not A202) );
 a8527a <=( A267  and  A266 );
 a8528a <=( a8527a  and  a8524a );
 a8531a <=( A199  and  A169 );
 a8534a <=( (not A201)  and  A200 );
 a8535a <=( a8534a  and  a8531a );
 a8538a <=( A232  and  (not A202) );
 a8541a <=( A301  and  A234 );
 a8542a <=( a8541a  and  a8538a );
 a8545a <=( A199  and  A169 );
 a8548a <=( (not A201)  and  A200 );
 a8549a <=( a8548a  and  a8545a );
 a8552a <=( A232  and  (not A202) );
 a8555a <=( A268  and  A234 );
 a8556a <=( a8555a  and  a8552a );
 a8559a <=( A199  and  A169 );
 a8562a <=( (not A201)  and  A200 );
 a8563a <=( a8562a  and  a8559a );
 a8566a <=( A233  and  (not A202) );
 a8569a <=( A301  and  A234 );
 a8570a <=( a8569a  and  a8566a );
 a8573a <=( A199  and  A169 );
 a8576a <=( (not A201)  and  A200 );
 a8577a <=( a8576a  and  a8573a );
 a8580a <=( A233  and  (not A202) );
 a8583a <=( A268  and  A234 );
 a8584a <=( a8583a  and  a8580a );
 a8587a <=( (not A199)  and  A169 );
 a8590a <=( (not A202)  and  (not A200) );
 a8591a <=( a8590a  and  a8587a );
 a8594a <=( A298  and  A235 );
 a8597a <=( A302  and  (not A299) );
 a8598a <=( a8597a  and  a8594a );
 a8601a <=( (not A199)  and  A169 );
 a8604a <=( (not A202)  and  (not A200) );
 a8605a <=( a8604a  and  a8601a );
 a8608a <=( (not A298)  and  A235 );
 a8611a <=( A302  and  A299 );
 a8612a <=( a8611a  and  a8608a );
 a8615a <=( (not A199)  and  A169 );
 a8618a <=( (not A202)  and  (not A200) );
 a8619a <=( a8618a  and  a8615a );
 a8622a <=( (not A265)  and  A235 );
 a8625a <=( A269  and  A266 );
 a8626a <=( a8625a  and  a8622a );
 a8629a <=( (not A199)  and  A169 );
 a8632a <=( (not A202)  and  (not A200) );
 a8633a <=( a8632a  and  a8629a );
 a8636a <=( A265  and  A235 );
 a8639a <=( A269  and  (not A266) );
 a8640a <=( a8639a  and  a8636a );
 a8643a <=( (not A199)  and  A169 );
 a8646a <=( (not A202)  and  (not A200) );
 a8647a <=( a8646a  and  a8643a );
 a8650a <=( A234  and  A232 );
 a8653a <=( A300  and  A299 );
 a8654a <=( a8653a  and  a8650a );
 a8657a <=( (not A199)  and  A169 );
 a8660a <=( (not A202)  and  (not A200) );
 a8661a <=( a8660a  and  a8657a );
 a8664a <=( A234  and  A232 );
 a8667a <=( A300  and  A298 );
 a8668a <=( a8667a  and  a8664a );
 a8671a <=( (not A199)  and  A169 );
 a8674a <=( (not A202)  and  (not A200) );
 a8675a <=( a8674a  and  a8671a );
 a8678a <=( A234  and  A232 );
 a8681a <=( A267  and  A265 );
 a8682a <=( a8681a  and  a8678a );
 a8685a <=( (not A199)  and  A169 );
 a8688a <=( (not A202)  and  (not A200) );
 a8689a <=( a8688a  and  a8685a );
 a8692a <=( A234  and  A232 );
 a8695a <=( A267  and  A266 );
 a8696a <=( a8695a  and  a8692a );
 a8699a <=( (not A199)  and  A169 );
 a8702a <=( (not A202)  and  (not A200) );
 a8703a <=( a8702a  and  a8699a );
 a8706a <=( A234  and  A233 );
 a8709a <=( A300  and  A299 );
 a8710a <=( a8709a  and  a8706a );
 a8713a <=( (not A199)  and  A169 );
 a8716a <=( (not A202)  and  (not A200) );
 a8717a <=( a8716a  and  a8713a );
 a8720a <=( A234  and  A233 );
 a8723a <=( A300  and  A298 );
 a8724a <=( a8723a  and  a8720a );
 a8727a <=( (not A199)  and  A169 );
 a8730a <=( (not A202)  and  (not A200) );
 a8731a <=( a8730a  and  a8727a );
 a8734a <=( A234  and  A233 );
 a8737a <=( A267  and  A265 );
 a8738a <=( a8737a  and  a8734a );
 a8741a <=( (not A199)  and  A169 );
 a8744a <=( (not A202)  and  (not A200) );
 a8745a <=( a8744a  and  a8741a );
 a8748a <=( A234  and  A233 );
 a8751a <=( A267  and  A266 );
 a8752a <=( a8751a  and  a8748a );
 a8755a <=( (not A199)  and  A169 );
 a8758a <=( (not A202)  and  (not A200) );
 a8759a <=( a8758a  and  a8755a );
 a8762a <=( A233  and  (not A232) );
 a8765a <=( A301  and  A236 );
 a8766a <=( a8765a  and  a8762a );
 a8769a <=( (not A199)  and  A169 );
 a8772a <=( (not A202)  and  (not A200) );
 a8773a <=( a8772a  and  a8769a );
 a8776a <=( A233  and  (not A232) );
 a8779a <=( A268  and  A236 );
 a8780a <=( a8779a  and  a8776a );
 a8783a <=( (not A199)  and  A169 );
 a8786a <=( (not A202)  and  (not A200) );
 a8787a <=( a8786a  and  a8783a );
 a8790a <=( (not A233)  and  A232 );
 a8793a <=( A301  and  A236 );
 a8794a <=( a8793a  and  a8790a );
 a8797a <=( (not A199)  and  A169 );
 a8800a <=( (not A202)  and  (not A200) );
 a8801a <=( a8800a  and  a8797a );
 a8804a <=( (not A233)  and  A232 );
 a8807a <=( A268  and  A236 );
 a8808a <=( a8807a  and  a8804a );
 a8811a <=( (not A167)  and  (not A169) );
 a8814a <=( A202  and  (not A166) );
 a8815a <=( a8814a  and  a8811a );
 a8818a <=( A298  and  A235 );
 a8821a <=( A302  and  (not A299) );
 a8822a <=( a8821a  and  a8818a );
 a8825a <=( (not A167)  and  (not A169) );
 a8828a <=( A202  and  (not A166) );
 a8829a <=( a8828a  and  a8825a );
 a8832a <=( (not A298)  and  A235 );
 a8835a <=( A302  and  A299 );
 a8836a <=( a8835a  and  a8832a );
 a8839a <=( (not A167)  and  (not A169) );
 a8842a <=( A202  and  (not A166) );
 a8843a <=( a8842a  and  a8839a );
 a8846a <=( (not A265)  and  A235 );
 a8849a <=( A269  and  A266 );
 a8850a <=( a8849a  and  a8846a );
 a8853a <=( (not A167)  and  (not A169) );
 a8856a <=( A202  and  (not A166) );
 a8857a <=( a8856a  and  a8853a );
 a8860a <=( A265  and  A235 );
 a8863a <=( A269  and  (not A266) );
 a8864a <=( a8863a  and  a8860a );
 a8867a <=( (not A167)  and  (not A169) );
 a8870a <=( A202  and  (not A166) );
 a8871a <=( a8870a  and  a8867a );
 a8874a <=( A234  and  A232 );
 a8877a <=( A300  and  A299 );
 a8878a <=( a8877a  and  a8874a );
 a8881a <=( (not A167)  and  (not A169) );
 a8884a <=( A202  and  (not A166) );
 a8885a <=( a8884a  and  a8881a );
 a8888a <=( A234  and  A232 );
 a8891a <=( A300  and  A298 );
 a8892a <=( a8891a  and  a8888a );
 a8895a <=( (not A167)  and  (not A169) );
 a8898a <=( A202  and  (not A166) );
 a8899a <=( a8898a  and  a8895a );
 a8902a <=( A234  and  A232 );
 a8905a <=( A267  and  A265 );
 a8906a <=( a8905a  and  a8902a );
 a8909a <=( (not A167)  and  (not A169) );
 a8912a <=( A202  and  (not A166) );
 a8913a <=( a8912a  and  a8909a );
 a8916a <=( A234  and  A232 );
 a8919a <=( A267  and  A266 );
 a8920a <=( a8919a  and  a8916a );
 a8923a <=( (not A167)  and  (not A169) );
 a8926a <=( A202  and  (not A166) );
 a8927a <=( a8926a  and  a8923a );
 a8930a <=( A234  and  A233 );
 a8933a <=( A300  and  A299 );
 a8934a <=( a8933a  and  a8930a );
 a8937a <=( (not A167)  and  (not A169) );
 a8940a <=( A202  and  (not A166) );
 a8941a <=( a8940a  and  a8937a );
 a8944a <=( A234  and  A233 );
 a8947a <=( A300  and  A298 );
 a8948a <=( a8947a  and  a8944a );
 a8951a <=( (not A167)  and  (not A169) );
 a8954a <=( A202  and  (not A166) );
 a8955a <=( a8954a  and  a8951a );
 a8958a <=( A234  and  A233 );
 a8961a <=( A267  and  A265 );
 a8962a <=( a8961a  and  a8958a );
 a8965a <=( (not A167)  and  (not A169) );
 a8968a <=( A202  and  (not A166) );
 a8969a <=( a8968a  and  a8965a );
 a8972a <=( A234  and  A233 );
 a8975a <=( A267  and  A266 );
 a8976a <=( a8975a  and  a8972a );
 a8979a <=( (not A167)  and  (not A169) );
 a8982a <=( A202  and  (not A166) );
 a8983a <=( a8982a  and  a8979a );
 a8986a <=( A233  and  (not A232) );
 a8989a <=( A301  and  A236 );
 a8990a <=( a8989a  and  a8986a );
 a8993a <=( (not A167)  and  (not A169) );
 a8996a <=( A202  and  (not A166) );
 a8997a <=( a8996a  and  a8993a );
 a9000a <=( A233  and  (not A232) );
 a9003a <=( A268  and  A236 );
 a9004a <=( a9003a  and  a9000a );
 a9007a <=( (not A167)  and  (not A169) );
 a9010a <=( A202  and  (not A166) );
 a9011a <=( a9010a  and  a9007a );
 a9014a <=( (not A233)  and  A232 );
 a9017a <=( A301  and  A236 );
 a9018a <=( a9017a  and  a9014a );
 a9021a <=( (not A167)  and  (not A169) );
 a9024a <=( A202  and  (not A166) );
 a9025a <=( a9024a  and  a9021a );
 a9028a <=( (not A233)  and  A232 );
 a9031a <=( A268  and  A236 );
 a9032a <=( a9031a  and  a9028a );
 a9035a <=( (not A167)  and  (not A169) );
 a9038a <=( A199  and  (not A166) );
 a9039a <=( a9038a  and  a9035a );
 a9042a <=( A235  and  A201 );
 a9045a <=( A300  and  A299 );
 a9046a <=( a9045a  and  a9042a );
 a9049a <=( (not A167)  and  (not A169) );
 a9052a <=( A199  and  (not A166) );
 a9053a <=( a9052a  and  a9049a );
 a9056a <=( A235  and  A201 );
 a9059a <=( A300  and  A298 );
 a9060a <=( a9059a  and  a9056a );
 a9063a <=( (not A167)  and  (not A169) );
 a9066a <=( A199  and  (not A166) );
 a9067a <=( a9066a  and  a9063a );
 a9070a <=( A235  and  A201 );
 a9073a <=( A267  and  A265 );
 a9074a <=( a9073a  and  a9070a );
 a9077a <=( (not A167)  and  (not A169) );
 a9080a <=( A199  and  (not A166) );
 a9081a <=( a9080a  and  a9077a );
 a9084a <=( A235  and  A201 );
 a9087a <=( A267  and  A266 );
 a9088a <=( a9087a  and  a9084a );
 a9091a <=( (not A167)  and  (not A169) );
 a9094a <=( A199  and  (not A166) );
 a9095a <=( a9094a  and  a9091a );
 a9098a <=( A232  and  A201 );
 a9101a <=( A301  and  A234 );
 a9102a <=( a9101a  and  a9098a );
 a9105a <=( (not A167)  and  (not A169) );
 a9108a <=( A199  and  (not A166) );
 a9109a <=( a9108a  and  a9105a );
 a9112a <=( A232  and  A201 );
 a9115a <=( A268  and  A234 );
 a9116a <=( a9115a  and  a9112a );
 a9119a <=( (not A167)  and  (not A169) );
 a9122a <=( A199  and  (not A166) );
 a9123a <=( a9122a  and  a9119a );
 a9126a <=( A233  and  A201 );
 a9129a <=( A301  and  A234 );
 a9130a <=( a9129a  and  a9126a );
 a9133a <=( (not A167)  and  (not A169) );
 a9136a <=( A199  and  (not A166) );
 a9137a <=( a9136a  and  a9133a );
 a9140a <=( A233  and  A201 );
 a9143a <=( A268  and  A234 );
 a9144a <=( a9143a  and  a9140a );
 a9147a <=( (not A167)  and  (not A169) );
 a9150a <=( A200  and  (not A166) );
 a9151a <=( a9150a  and  a9147a );
 a9154a <=( A235  and  A201 );
 a9157a <=( A300  and  A299 );
 a9158a <=( a9157a  and  a9154a );
 a9161a <=( (not A167)  and  (not A169) );
 a9164a <=( A200  and  (not A166) );
 a9165a <=( a9164a  and  a9161a );
 a9168a <=( A235  and  A201 );
 a9171a <=( A300  and  A298 );
 a9172a <=( a9171a  and  a9168a );
 a9175a <=( (not A167)  and  (not A169) );
 a9178a <=( A200  and  (not A166) );
 a9179a <=( a9178a  and  a9175a );
 a9182a <=( A235  and  A201 );
 a9185a <=( A267  and  A265 );
 a9186a <=( a9185a  and  a9182a );
 a9189a <=( (not A167)  and  (not A169) );
 a9192a <=( A200  and  (not A166) );
 a9193a <=( a9192a  and  a9189a );
 a9196a <=( A235  and  A201 );
 a9199a <=( A267  and  A266 );
 a9200a <=( a9199a  and  a9196a );
 a9203a <=( (not A167)  and  (not A169) );
 a9206a <=( A200  and  (not A166) );
 a9207a <=( a9206a  and  a9203a );
 a9210a <=( A232  and  A201 );
 a9213a <=( A301  and  A234 );
 a9214a <=( a9213a  and  a9210a );
 a9217a <=( (not A167)  and  (not A169) );
 a9220a <=( A200  and  (not A166) );
 a9221a <=( a9220a  and  a9217a );
 a9224a <=( A232  and  A201 );
 a9227a <=( A268  and  A234 );
 a9228a <=( a9227a  and  a9224a );
 a9231a <=( (not A167)  and  (not A169) );
 a9234a <=( A200  and  (not A166) );
 a9235a <=( a9234a  and  a9231a );
 a9238a <=( A233  and  A201 );
 a9241a <=( A301  and  A234 );
 a9242a <=( a9241a  and  a9238a );
 a9245a <=( (not A167)  and  (not A169) );
 a9248a <=( A200  and  (not A166) );
 a9249a <=( a9248a  and  a9245a );
 a9252a <=( A233  and  A201 );
 a9255a <=( A268  and  A234 );
 a9256a <=( a9255a  and  a9252a );
 a9259a <=( (not A167)  and  (not A169) );
 a9262a <=( (not A199)  and  (not A166) );
 a9263a <=( a9262a  and  a9259a );
 a9266a <=( A203  and  A200 );
 a9269a <=( A301  and  A235 );
 a9270a <=( a9269a  and  a9266a );
 a9273a <=( (not A167)  and  (not A169) );
 a9276a <=( (not A199)  and  (not A166) );
 a9277a <=( a9276a  and  a9273a );
 a9280a <=( A203  and  A200 );
 a9283a <=( A268  and  A235 );
 a9284a <=( a9283a  and  a9280a );
 a9287a <=( (not A167)  and  (not A169) );
 a9290a <=( A199  and  (not A166) );
 a9291a <=( a9290a  and  a9287a );
 a9294a <=( A203  and  (not A200) );
 a9297a <=( A301  and  A235 );
 a9298a <=( a9297a  and  a9294a );
 a9301a <=( (not A167)  and  (not A169) );
 a9304a <=( A199  and  (not A166) );
 a9305a <=( a9304a  and  a9301a );
 a9308a <=( A203  and  (not A200) );
 a9311a <=( A268  and  A235 );
 a9312a <=( a9311a  and  a9308a );
 a9315a <=( (not A168)  and  (not A169) );
 a9318a <=( A166  and  A167 );
 a9319a <=( a9318a  and  a9315a );
 a9322a <=( A235  and  A202 );
 a9325a <=( A300  and  A299 );
 a9326a <=( a9325a  and  a9322a );
 a9329a <=( (not A168)  and  (not A169) );
 a9332a <=( A166  and  A167 );
 a9333a <=( a9332a  and  a9329a );
 a9336a <=( A235  and  A202 );
 a9339a <=( A300  and  A298 );
 a9340a <=( a9339a  and  a9336a );
 a9343a <=( (not A168)  and  (not A169) );
 a9346a <=( A166  and  A167 );
 a9347a <=( a9346a  and  a9343a );
 a9350a <=( A235  and  A202 );
 a9353a <=( A267  and  A265 );
 a9354a <=( a9353a  and  a9350a );
 a9357a <=( (not A168)  and  (not A169) );
 a9360a <=( A166  and  A167 );
 a9361a <=( a9360a  and  a9357a );
 a9364a <=( A235  and  A202 );
 a9367a <=( A267  and  A266 );
 a9368a <=( a9367a  and  a9364a );
 a9371a <=( (not A168)  and  (not A169) );
 a9374a <=( A166  and  A167 );
 a9375a <=( a9374a  and  a9371a );
 a9378a <=( A232  and  A202 );
 a9381a <=( A301  and  A234 );
 a9382a <=( a9381a  and  a9378a );
 a9385a <=( (not A168)  and  (not A169) );
 a9388a <=( A166  and  A167 );
 a9389a <=( a9388a  and  a9385a );
 a9392a <=( A232  and  A202 );
 a9395a <=( A268  and  A234 );
 a9396a <=( a9395a  and  a9392a );
 a9399a <=( (not A168)  and  (not A169) );
 a9402a <=( A166  and  A167 );
 a9403a <=( a9402a  and  a9399a );
 a9406a <=( A233  and  A202 );
 a9409a <=( A301  and  A234 );
 a9410a <=( a9409a  and  a9406a );
 a9413a <=( (not A168)  and  (not A169) );
 a9416a <=( A166  and  A167 );
 a9417a <=( a9416a  and  a9413a );
 a9420a <=( A233  and  A202 );
 a9423a <=( A268  and  A234 );
 a9424a <=( a9423a  and  a9420a );
 a9427a <=( (not A168)  and  (not A169) );
 a9430a <=( A166  and  A167 );
 a9431a <=( a9430a  and  a9427a );
 a9434a <=( A201  and  A199 );
 a9437a <=( A301  and  A235 );
 a9438a <=( a9437a  and  a9434a );
 a9441a <=( (not A168)  and  (not A169) );
 a9444a <=( A166  and  A167 );
 a9445a <=( a9444a  and  a9441a );
 a9448a <=( A201  and  A199 );
 a9451a <=( A268  and  A235 );
 a9452a <=( a9451a  and  a9448a );
 a9455a <=( (not A168)  and  (not A169) );
 a9458a <=( A166  and  A167 );
 a9459a <=( a9458a  and  a9455a );
 a9462a <=( A201  and  A200 );
 a9465a <=( A301  and  A235 );
 a9466a <=( a9465a  and  a9462a );
 a9469a <=( (not A168)  and  (not A169) );
 a9472a <=( A166  and  A167 );
 a9473a <=( a9472a  and  a9469a );
 a9476a <=( A201  and  A200 );
 a9479a <=( A268  and  A235 );
 a9480a <=( a9479a  and  a9476a );
 a9483a <=( (not A169)  and  (not A170) );
 a9486a <=( A202  and  (not A168) );
 a9487a <=( a9486a  and  a9483a );
 a9490a <=( A298  and  A235 );
 a9493a <=( A302  and  (not A299) );
 a9494a <=( a9493a  and  a9490a );
 a9497a <=( (not A169)  and  (not A170) );
 a9500a <=( A202  and  (not A168) );
 a9501a <=( a9500a  and  a9497a );
 a9504a <=( (not A298)  and  A235 );
 a9507a <=( A302  and  A299 );
 a9508a <=( a9507a  and  a9504a );
 a9511a <=( (not A169)  and  (not A170) );
 a9514a <=( A202  and  (not A168) );
 a9515a <=( a9514a  and  a9511a );
 a9518a <=( (not A265)  and  A235 );
 a9521a <=( A269  and  A266 );
 a9522a <=( a9521a  and  a9518a );
 a9525a <=( (not A169)  and  (not A170) );
 a9528a <=( A202  and  (not A168) );
 a9529a <=( a9528a  and  a9525a );
 a9532a <=( A265  and  A235 );
 a9535a <=( A269  and  (not A266) );
 a9536a <=( a9535a  and  a9532a );
 a9539a <=( (not A169)  and  (not A170) );
 a9542a <=( A202  and  (not A168) );
 a9543a <=( a9542a  and  a9539a );
 a9546a <=( A234  and  A232 );
 a9549a <=( A300  and  A299 );
 a9550a <=( a9549a  and  a9546a );
 a9553a <=( (not A169)  and  (not A170) );
 a9556a <=( A202  and  (not A168) );
 a9557a <=( a9556a  and  a9553a );
 a9560a <=( A234  and  A232 );
 a9563a <=( A300  and  A298 );
 a9564a <=( a9563a  and  a9560a );
 a9567a <=( (not A169)  and  (not A170) );
 a9570a <=( A202  and  (not A168) );
 a9571a <=( a9570a  and  a9567a );
 a9574a <=( A234  and  A232 );
 a9577a <=( A267  and  A265 );
 a9578a <=( a9577a  and  a9574a );
 a9581a <=( (not A169)  and  (not A170) );
 a9584a <=( A202  and  (not A168) );
 a9585a <=( a9584a  and  a9581a );
 a9588a <=( A234  and  A232 );
 a9591a <=( A267  and  A266 );
 a9592a <=( a9591a  and  a9588a );
 a9595a <=( (not A169)  and  (not A170) );
 a9598a <=( A202  and  (not A168) );
 a9599a <=( a9598a  and  a9595a );
 a9602a <=( A234  and  A233 );
 a9605a <=( A300  and  A299 );
 a9606a <=( a9605a  and  a9602a );
 a9609a <=( (not A169)  and  (not A170) );
 a9612a <=( A202  and  (not A168) );
 a9613a <=( a9612a  and  a9609a );
 a9616a <=( A234  and  A233 );
 a9619a <=( A300  and  A298 );
 a9620a <=( a9619a  and  a9616a );
 a9623a <=( (not A169)  and  (not A170) );
 a9626a <=( A202  and  (not A168) );
 a9627a <=( a9626a  and  a9623a );
 a9630a <=( A234  and  A233 );
 a9633a <=( A267  and  A265 );
 a9634a <=( a9633a  and  a9630a );
 a9637a <=( (not A169)  and  (not A170) );
 a9640a <=( A202  and  (not A168) );
 a9641a <=( a9640a  and  a9637a );
 a9644a <=( A234  and  A233 );
 a9647a <=( A267  and  A266 );
 a9648a <=( a9647a  and  a9644a );
 a9651a <=( (not A169)  and  (not A170) );
 a9654a <=( A202  and  (not A168) );
 a9655a <=( a9654a  and  a9651a );
 a9658a <=( A233  and  (not A232) );
 a9661a <=( A301  and  A236 );
 a9662a <=( a9661a  and  a9658a );
 a9665a <=( (not A169)  and  (not A170) );
 a9668a <=( A202  and  (not A168) );
 a9669a <=( a9668a  and  a9665a );
 a9672a <=( A233  and  (not A232) );
 a9675a <=( A268  and  A236 );
 a9676a <=( a9675a  and  a9672a );
 a9679a <=( (not A169)  and  (not A170) );
 a9682a <=( A202  and  (not A168) );
 a9683a <=( a9682a  and  a9679a );
 a9686a <=( (not A233)  and  A232 );
 a9689a <=( A301  and  A236 );
 a9690a <=( a9689a  and  a9686a );
 a9693a <=( (not A169)  and  (not A170) );
 a9696a <=( A202  and  (not A168) );
 a9697a <=( a9696a  and  a9693a );
 a9700a <=( (not A233)  and  A232 );
 a9703a <=( A268  and  A236 );
 a9704a <=( a9703a  and  a9700a );
 a9707a <=( (not A169)  and  (not A170) );
 a9710a <=( A199  and  (not A168) );
 a9711a <=( a9710a  and  a9707a );
 a9714a <=( A235  and  A201 );
 a9717a <=( A300  and  A299 );
 a9718a <=( a9717a  and  a9714a );
 a9721a <=( (not A169)  and  (not A170) );
 a9724a <=( A199  and  (not A168) );
 a9725a <=( a9724a  and  a9721a );
 a9728a <=( A235  and  A201 );
 a9731a <=( A300  and  A298 );
 a9732a <=( a9731a  and  a9728a );
 a9735a <=( (not A169)  and  (not A170) );
 a9738a <=( A199  and  (not A168) );
 a9739a <=( a9738a  and  a9735a );
 a9742a <=( A235  and  A201 );
 a9745a <=( A267  and  A265 );
 a9746a <=( a9745a  and  a9742a );
 a9749a <=( (not A169)  and  (not A170) );
 a9752a <=( A199  and  (not A168) );
 a9753a <=( a9752a  and  a9749a );
 a9756a <=( A235  and  A201 );
 a9759a <=( A267  and  A266 );
 a9760a <=( a9759a  and  a9756a );
 a9763a <=( (not A169)  and  (not A170) );
 a9766a <=( A199  and  (not A168) );
 a9767a <=( a9766a  and  a9763a );
 a9770a <=( A232  and  A201 );
 a9773a <=( A301  and  A234 );
 a9774a <=( a9773a  and  a9770a );
 a9777a <=( (not A169)  and  (not A170) );
 a9780a <=( A199  and  (not A168) );
 a9781a <=( a9780a  and  a9777a );
 a9784a <=( A232  and  A201 );
 a9787a <=( A268  and  A234 );
 a9788a <=( a9787a  and  a9784a );
 a9791a <=( (not A169)  and  (not A170) );
 a9794a <=( A199  and  (not A168) );
 a9795a <=( a9794a  and  a9791a );
 a9798a <=( A233  and  A201 );
 a9801a <=( A301  and  A234 );
 a9802a <=( a9801a  and  a9798a );
 a9805a <=( (not A169)  and  (not A170) );
 a9808a <=( A199  and  (not A168) );
 a9809a <=( a9808a  and  a9805a );
 a9812a <=( A233  and  A201 );
 a9815a <=( A268  and  A234 );
 a9816a <=( a9815a  and  a9812a );
 a9819a <=( (not A169)  and  (not A170) );
 a9822a <=( A200  and  (not A168) );
 a9823a <=( a9822a  and  a9819a );
 a9826a <=( A235  and  A201 );
 a9829a <=( A300  and  A299 );
 a9830a <=( a9829a  and  a9826a );
 a9833a <=( (not A169)  and  (not A170) );
 a9836a <=( A200  and  (not A168) );
 a9837a <=( a9836a  and  a9833a );
 a9840a <=( A235  and  A201 );
 a9843a <=( A300  and  A298 );
 a9844a <=( a9843a  and  a9840a );
 a9847a <=( (not A169)  and  (not A170) );
 a9850a <=( A200  and  (not A168) );
 a9851a <=( a9850a  and  a9847a );
 a9854a <=( A235  and  A201 );
 a9857a <=( A267  and  A265 );
 a9858a <=( a9857a  and  a9854a );
 a9861a <=( (not A169)  and  (not A170) );
 a9864a <=( A200  and  (not A168) );
 a9865a <=( a9864a  and  a9861a );
 a9868a <=( A235  and  A201 );
 a9871a <=( A267  and  A266 );
 a9872a <=( a9871a  and  a9868a );
 a9875a <=( (not A169)  and  (not A170) );
 a9878a <=( A200  and  (not A168) );
 a9879a <=( a9878a  and  a9875a );
 a9882a <=( A232  and  A201 );
 a9885a <=( A301  and  A234 );
 a9886a <=( a9885a  and  a9882a );
 a9889a <=( (not A169)  and  (not A170) );
 a9892a <=( A200  and  (not A168) );
 a9893a <=( a9892a  and  a9889a );
 a9896a <=( A232  and  A201 );
 a9899a <=( A268  and  A234 );
 a9900a <=( a9899a  and  a9896a );
 a9903a <=( (not A169)  and  (not A170) );
 a9906a <=( A200  and  (not A168) );
 a9907a <=( a9906a  and  a9903a );
 a9910a <=( A233  and  A201 );
 a9913a <=( A301  and  A234 );
 a9914a <=( a9913a  and  a9910a );
 a9917a <=( (not A169)  and  (not A170) );
 a9920a <=( A200  and  (not A168) );
 a9921a <=( a9920a  and  a9917a );
 a9924a <=( A233  and  A201 );
 a9927a <=( A268  and  A234 );
 a9928a <=( a9927a  and  a9924a );
 a9931a <=( (not A169)  and  (not A170) );
 a9934a <=( (not A199)  and  (not A168) );
 a9935a <=( a9934a  and  a9931a );
 a9938a <=( A203  and  A200 );
 a9941a <=( A301  and  A235 );
 a9942a <=( a9941a  and  a9938a );
 a9945a <=( (not A169)  and  (not A170) );
 a9948a <=( (not A199)  and  (not A168) );
 a9949a <=( a9948a  and  a9945a );
 a9952a <=( A203  and  A200 );
 a9955a <=( A268  and  A235 );
 a9956a <=( a9955a  and  a9952a );
 a9959a <=( (not A169)  and  (not A170) );
 a9962a <=( A199  and  (not A168) );
 a9963a <=( a9962a  and  a9959a );
 a9966a <=( A203  and  (not A200) );
 a9969a <=( A301  and  A235 );
 a9970a <=( a9969a  and  a9966a );
 a9973a <=( (not A169)  and  (not A170) );
 a9976a <=( A199  and  (not A168) );
 a9977a <=( a9976a  and  a9973a );
 a9980a <=( A203  and  (not A200) );
 a9983a <=( A268  and  A235 );
 a9984a <=( a9983a  and  a9980a );
 a9987a <=( A166  and  A168 );
 a9990a <=( (not A202)  and  (not A201) );
 a9991a <=( a9990a  and  a9987a );
 a9994a <=( A235  and  (not A203) );
 a9998a <=( A302  and  (not A299) );
 a9999a <=( A298  and  a9998a );
 a10000a <=( a9999a  and  a9994a );
 a10003a <=( A166  and  A168 );
 a10006a <=( (not A202)  and  (not A201) );
 a10007a <=( a10006a  and  a10003a );
 a10010a <=( A235  and  (not A203) );
 a10014a <=( A302  and  A299 );
 a10015a <=( (not A298)  and  a10014a );
 a10016a <=( a10015a  and  a10010a );
 a10019a <=( A166  and  A168 );
 a10022a <=( (not A202)  and  (not A201) );
 a10023a <=( a10022a  and  a10019a );
 a10026a <=( A235  and  (not A203) );
 a10030a <=( A269  and  A266 );
 a10031a <=( (not A265)  and  a10030a );
 a10032a <=( a10031a  and  a10026a );
 a10035a <=( A166  and  A168 );
 a10038a <=( (not A202)  and  (not A201) );
 a10039a <=( a10038a  and  a10035a );
 a10042a <=( A235  and  (not A203) );
 a10046a <=( A269  and  (not A266) );
 a10047a <=( A265  and  a10046a );
 a10048a <=( a10047a  and  a10042a );
 a10051a <=( A166  and  A168 );
 a10054a <=( (not A202)  and  (not A201) );
 a10055a <=( a10054a  and  a10051a );
 a10058a <=( A232  and  (not A203) );
 a10062a <=( A300  and  A299 );
 a10063a <=( A234  and  a10062a );
 a10064a <=( a10063a  and  a10058a );
 a10067a <=( A166  and  A168 );
 a10070a <=( (not A202)  and  (not A201) );
 a10071a <=( a10070a  and  a10067a );
 a10074a <=( A232  and  (not A203) );
 a10078a <=( A300  and  A298 );
 a10079a <=( A234  and  a10078a );
 a10080a <=( a10079a  and  a10074a );
 a10083a <=( A166  and  A168 );
 a10086a <=( (not A202)  and  (not A201) );
 a10087a <=( a10086a  and  a10083a );
 a10090a <=( A232  and  (not A203) );
 a10094a <=( A267  and  A265 );
 a10095a <=( A234  and  a10094a );
 a10096a <=( a10095a  and  a10090a );
 a10099a <=( A166  and  A168 );
 a10102a <=( (not A202)  and  (not A201) );
 a10103a <=( a10102a  and  a10099a );
 a10106a <=( A232  and  (not A203) );
 a10110a <=( A267  and  A266 );
 a10111a <=( A234  and  a10110a );
 a10112a <=( a10111a  and  a10106a );
 a10115a <=( A166  and  A168 );
 a10118a <=( (not A202)  and  (not A201) );
 a10119a <=( a10118a  and  a10115a );
 a10122a <=( A233  and  (not A203) );
 a10126a <=( A300  and  A299 );
 a10127a <=( A234  and  a10126a );
 a10128a <=( a10127a  and  a10122a );
 a10131a <=( A166  and  A168 );
 a10134a <=( (not A202)  and  (not A201) );
 a10135a <=( a10134a  and  a10131a );
 a10138a <=( A233  and  (not A203) );
 a10142a <=( A300  and  A298 );
 a10143a <=( A234  and  a10142a );
 a10144a <=( a10143a  and  a10138a );
 a10147a <=( A166  and  A168 );
 a10150a <=( (not A202)  and  (not A201) );
 a10151a <=( a10150a  and  a10147a );
 a10154a <=( A233  and  (not A203) );
 a10158a <=( A267  and  A265 );
 a10159a <=( A234  and  a10158a );
 a10160a <=( a10159a  and  a10154a );
 a10163a <=( A166  and  A168 );
 a10166a <=( (not A202)  and  (not A201) );
 a10167a <=( a10166a  and  a10163a );
 a10170a <=( A233  and  (not A203) );
 a10174a <=( A267  and  A266 );
 a10175a <=( A234  and  a10174a );
 a10176a <=( a10175a  and  a10170a );
 a10179a <=( A166  and  A168 );
 a10182a <=( (not A202)  and  (not A201) );
 a10183a <=( a10182a  and  a10179a );
 a10186a <=( (not A232)  and  (not A203) );
 a10190a <=( A301  and  A236 );
 a10191a <=( A233  and  a10190a );
 a10192a <=( a10191a  and  a10186a );
 a10195a <=( A166  and  A168 );
 a10198a <=( (not A202)  and  (not A201) );
 a10199a <=( a10198a  and  a10195a );
 a10202a <=( (not A232)  and  (not A203) );
 a10206a <=( A268  and  A236 );
 a10207a <=( A233  and  a10206a );
 a10208a <=( a10207a  and  a10202a );
 a10211a <=( A166  and  A168 );
 a10214a <=( (not A202)  and  (not A201) );
 a10215a <=( a10214a  and  a10211a );
 a10218a <=( A232  and  (not A203) );
 a10222a <=( A301  and  A236 );
 a10223a <=( (not A233)  and  a10222a );
 a10224a <=( a10223a  and  a10218a );
 a10227a <=( A166  and  A168 );
 a10230a <=( (not A202)  and  (not A201) );
 a10231a <=( a10230a  and  a10227a );
 a10234a <=( A232  and  (not A203) );
 a10238a <=( A268  and  A236 );
 a10239a <=( (not A233)  and  a10238a );
 a10240a <=( a10239a  and  a10234a );
 a10243a <=( A166  and  A168 );
 a10246a <=( A200  and  A199 );
 a10247a <=( a10246a  and  a10243a );
 a10250a <=( (not A202)  and  (not A201) );
 a10254a <=( A300  and  A299 );
 a10255a <=( A235  and  a10254a );
 a10256a <=( a10255a  and  a10250a );
 a10259a <=( A166  and  A168 );
 a10262a <=( A200  and  A199 );
 a10263a <=( a10262a  and  a10259a );
 a10266a <=( (not A202)  and  (not A201) );
 a10270a <=( A300  and  A298 );
 a10271a <=( A235  and  a10270a );
 a10272a <=( a10271a  and  a10266a );
 a10275a <=( A166  and  A168 );
 a10278a <=( A200  and  A199 );
 a10279a <=( a10278a  and  a10275a );
 a10282a <=( (not A202)  and  (not A201) );
 a10286a <=( A267  and  A265 );
 a10287a <=( A235  and  a10286a );
 a10288a <=( a10287a  and  a10282a );
 a10291a <=( A166  and  A168 );
 a10294a <=( A200  and  A199 );
 a10295a <=( a10294a  and  a10291a );
 a10298a <=( (not A202)  and  (not A201) );
 a10302a <=( A267  and  A266 );
 a10303a <=( A235  and  a10302a );
 a10304a <=( a10303a  and  a10298a );
 a10307a <=( A166  and  A168 );
 a10310a <=( A200  and  A199 );
 a10311a <=( a10310a  and  a10307a );
 a10314a <=( (not A202)  and  (not A201) );
 a10318a <=( A301  and  A234 );
 a10319a <=( A232  and  a10318a );
 a10320a <=( a10319a  and  a10314a );
 a10323a <=( A166  and  A168 );
 a10326a <=( A200  and  A199 );
 a10327a <=( a10326a  and  a10323a );
 a10330a <=( (not A202)  and  (not A201) );
 a10334a <=( A268  and  A234 );
 a10335a <=( A232  and  a10334a );
 a10336a <=( a10335a  and  a10330a );
 a10339a <=( A166  and  A168 );
 a10342a <=( A200  and  A199 );
 a10343a <=( a10342a  and  a10339a );
 a10346a <=( (not A202)  and  (not A201) );
 a10350a <=( A301  and  A234 );
 a10351a <=( A233  and  a10350a );
 a10352a <=( a10351a  and  a10346a );
 a10355a <=( A166  and  A168 );
 a10358a <=( A200  and  A199 );
 a10359a <=( a10358a  and  a10355a );
 a10362a <=( (not A202)  and  (not A201) );
 a10366a <=( A268  and  A234 );
 a10367a <=( A233  and  a10366a );
 a10368a <=( a10367a  and  a10362a );
 a10371a <=( A166  and  A168 );
 a10374a <=( (not A200)  and  (not A199) );
 a10375a <=( a10374a  and  a10371a );
 a10378a <=( A235  and  (not A202) );
 a10382a <=( A302  and  (not A299) );
 a10383a <=( A298  and  a10382a );
 a10384a <=( a10383a  and  a10378a );
 a10387a <=( A166  and  A168 );
 a10390a <=( (not A200)  and  (not A199) );
 a10391a <=( a10390a  and  a10387a );
 a10394a <=( A235  and  (not A202) );
 a10398a <=( A302  and  A299 );
 a10399a <=( (not A298)  and  a10398a );
 a10400a <=( a10399a  and  a10394a );
 a10403a <=( A166  and  A168 );
 a10406a <=( (not A200)  and  (not A199) );
 a10407a <=( a10406a  and  a10403a );
 a10410a <=( A235  and  (not A202) );
 a10414a <=( A269  and  A266 );
 a10415a <=( (not A265)  and  a10414a );
 a10416a <=( a10415a  and  a10410a );
 a10419a <=( A166  and  A168 );
 a10422a <=( (not A200)  and  (not A199) );
 a10423a <=( a10422a  and  a10419a );
 a10426a <=( A235  and  (not A202) );
 a10430a <=( A269  and  (not A266) );
 a10431a <=( A265  and  a10430a );
 a10432a <=( a10431a  and  a10426a );
 a10435a <=( A166  and  A168 );
 a10438a <=( (not A200)  and  (not A199) );
 a10439a <=( a10438a  and  a10435a );
 a10442a <=( A232  and  (not A202) );
 a10446a <=( A300  and  A299 );
 a10447a <=( A234  and  a10446a );
 a10448a <=( a10447a  and  a10442a );
 a10451a <=( A166  and  A168 );
 a10454a <=( (not A200)  and  (not A199) );
 a10455a <=( a10454a  and  a10451a );
 a10458a <=( A232  and  (not A202) );
 a10462a <=( A300  and  A298 );
 a10463a <=( A234  and  a10462a );
 a10464a <=( a10463a  and  a10458a );
 a10467a <=( A166  and  A168 );
 a10470a <=( (not A200)  and  (not A199) );
 a10471a <=( a10470a  and  a10467a );
 a10474a <=( A232  and  (not A202) );
 a10478a <=( A267  and  A265 );
 a10479a <=( A234  and  a10478a );
 a10480a <=( a10479a  and  a10474a );
 a10483a <=( A166  and  A168 );
 a10486a <=( (not A200)  and  (not A199) );
 a10487a <=( a10486a  and  a10483a );
 a10490a <=( A232  and  (not A202) );
 a10494a <=( A267  and  A266 );
 a10495a <=( A234  and  a10494a );
 a10496a <=( a10495a  and  a10490a );
 a10499a <=( A166  and  A168 );
 a10502a <=( (not A200)  and  (not A199) );
 a10503a <=( a10502a  and  a10499a );
 a10506a <=( A233  and  (not A202) );
 a10510a <=( A300  and  A299 );
 a10511a <=( A234  and  a10510a );
 a10512a <=( a10511a  and  a10506a );
 a10515a <=( A166  and  A168 );
 a10518a <=( (not A200)  and  (not A199) );
 a10519a <=( a10518a  and  a10515a );
 a10522a <=( A233  and  (not A202) );
 a10526a <=( A300  and  A298 );
 a10527a <=( A234  and  a10526a );
 a10528a <=( a10527a  and  a10522a );
 a10531a <=( A166  and  A168 );
 a10534a <=( (not A200)  and  (not A199) );
 a10535a <=( a10534a  and  a10531a );
 a10538a <=( A233  and  (not A202) );
 a10542a <=( A267  and  A265 );
 a10543a <=( A234  and  a10542a );
 a10544a <=( a10543a  and  a10538a );
 a10547a <=( A166  and  A168 );
 a10550a <=( (not A200)  and  (not A199) );
 a10551a <=( a10550a  and  a10547a );
 a10554a <=( A233  and  (not A202) );
 a10558a <=( A267  and  A266 );
 a10559a <=( A234  and  a10558a );
 a10560a <=( a10559a  and  a10554a );
 a10563a <=( A166  and  A168 );
 a10566a <=( (not A200)  and  (not A199) );
 a10567a <=( a10566a  and  a10563a );
 a10570a <=( (not A232)  and  (not A202) );
 a10574a <=( A301  and  A236 );
 a10575a <=( A233  and  a10574a );
 a10576a <=( a10575a  and  a10570a );
 a10579a <=( A166  and  A168 );
 a10582a <=( (not A200)  and  (not A199) );
 a10583a <=( a10582a  and  a10579a );
 a10586a <=( (not A232)  and  (not A202) );
 a10590a <=( A268  and  A236 );
 a10591a <=( A233  and  a10590a );
 a10592a <=( a10591a  and  a10586a );
 a10595a <=( A166  and  A168 );
 a10598a <=( (not A200)  and  (not A199) );
 a10599a <=( a10598a  and  a10595a );
 a10602a <=( A232  and  (not A202) );
 a10606a <=( A301  and  A236 );
 a10607a <=( (not A233)  and  a10606a );
 a10608a <=( a10607a  and  a10602a );
 a10611a <=( A166  and  A168 );
 a10614a <=( (not A200)  and  (not A199) );
 a10615a <=( a10614a  and  a10611a );
 a10618a <=( A232  and  (not A202) );
 a10622a <=( A268  and  A236 );
 a10623a <=( (not A233)  and  a10622a );
 a10624a <=( a10623a  and  a10618a );
 a10627a <=( A167  and  A168 );
 a10630a <=( (not A202)  and  (not A201) );
 a10631a <=( a10630a  and  a10627a );
 a10634a <=( A235  and  (not A203) );
 a10638a <=( A302  and  (not A299) );
 a10639a <=( A298  and  a10638a );
 a10640a <=( a10639a  and  a10634a );
 a10643a <=( A167  and  A168 );
 a10646a <=( (not A202)  and  (not A201) );
 a10647a <=( a10646a  and  a10643a );
 a10650a <=( A235  and  (not A203) );
 a10654a <=( A302  and  A299 );
 a10655a <=( (not A298)  and  a10654a );
 a10656a <=( a10655a  and  a10650a );
 a10659a <=( A167  and  A168 );
 a10662a <=( (not A202)  and  (not A201) );
 a10663a <=( a10662a  and  a10659a );
 a10666a <=( A235  and  (not A203) );
 a10670a <=( A269  and  A266 );
 a10671a <=( (not A265)  and  a10670a );
 a10672a <=( a10671a  and  a10666a );
 a10675a <=( A167  and  A168 );
 a10678a <=( (not A202)  and  (not A201) );
 a10679a <=( a10678a  and  a10675a );
 a10682a <=( A235  and  (not A203) );
 a10686a <=( A269  and  (not A266) );
 a10687a <=( A265  and  a10686a );
 a10688a <=( a10687a  and  a10682a );
 a10691a <=( A167  and  A168 );
 a10694a <=( (not A202)  and  (not A201) );
 a10695a <=( a10694a  and  a10691a );
 a10698a <=( A232  and  (not A203) );
 a10702a <=( A300  and  A299 );
 a10703a <=( A234  and  a10702a );
 a10704a <=( a10703a  and  a10698a );
 a10707a <=( A167  and  A168 );
 a10710a <=( (not A202)  and  (not A201) );
 a10711a <=( a10710a  and  a10707a );
 a10714a <=( A232  and  (not A203) );
 a10718a <=( A300  and  A298 );
 a10719a <=( A234  and  a10718a );
 a10720a <=( a10719a  and  a10714a );
 a10723a <=( A167  and  A168 );
 a10726a <=( (not A202)  and  (not A201) );
 a10727a <=( a10726a  and  a10723a );
 a10730a <=( A232  and  (not A203) );
 a10734a <=( A267  and  A265 );
 a10735a <=( A234  and  a10734a );
 a10736a <=( a10735a  and  a10730a );
 a10739a <=( A167  and  A168 );
 a10742a <=( (not A202)  and  (not A201) );
 a10743a <=( a10742a  and  a10739a );
 a10746a <=( A232  and  (not A203) );
 a10750a <=( A267  and  A266 );
 a10751a <=( A234  and  a10750a );
 a10752a <=( a10751a  and  a10746a );
 a10755a <=( A167  and  A168 );
 a10758a <=( (not A202)  and  (not A201) );
 a10759a <=( a10758a  and  a10755a );
 a10762a <=( A233  and  (not A203) );
 a10766a <=( A300  and  A299 );
 a10767a <=( A234  and  a10766a );
 a10768a <=( a10767a  and  a10762a );
 a10771a <=( A167  and  A168 );
 a10774a <=( (not A202)  and  (not A201) );
 a10775a <=( a10774a  and  a10771a );
 a10778a <=( A233  and  (not A203) );
 a10782a <=( A300  and  A298 );
 a10783a <=( A234  and  a10782a );
 a10784a <=( a10783a  and  a10778a );
 a10787a <=( A167  and  A168 );
 a10790a <=( (not A202)  and  (not A201) );
 a10791a <=( a10790a  and  a10787a );
 a10794a <=( A233  and  (not A203) );
 a10798a <=( A267  and  A265 );
 a10799a <=( A234  and  a10798a );
 a10800a <=( a10799a  and  a10794a );
 a10803a <=( A167  and  A168 );
 a10806a <=( (not A202)  and  (not A201) );
 a10807a <=( a10806a  and  a10803a );
 a10810a <=( A233  and  (not A203) );
 a10814a <=( A267  and  A266 );
 a10815a <=( A234  and  a10814a );
 a10816a <=( a10815a  and  a10810a );
 a10819a <=( A167  and  A168 );
 a10822a <=( (not A202)  and  (not A201) );
 a10823a <=( a10822a  and  a10819a );
 a10826a <=( (not A232)  and  (not A203) );
 a10830a <=( A301  and  A236 );
 a10831a <=( A233  and  a10830a );
 a10832a <=( a10831a  and  a10826a );
 a10835a <=( A167  and  A168 );
 a10838a <=( (not A202)  and  (not A201) );
 a10839a <=( a10838a  and  a10835a );
 a10842a <=( (not A232)  and  (not A203) );
 a10846a <=( A268  and  A236 );
 a10847a <=( A233  and  a10846a );
 a10848a <=( a10847a  and  a10842a );
 a10851a <=( A167  and  A168 );
 a10854a <=( (not A202)  and  (not A201) );
 a10855a <=( a10854a  and  a10851a );
 a10858a <=( A232  and  (not A203) );
 a10862a <=( A301  and  A236 );
 a10863a <=( (not A233)  and  a10862a );
 a10864a <=( a10863a  and  a10858a );
 a10867a <=( A167  and  A168 );
 a10870a <=( (not A202)  and  (not A201) );
 a10871a <=( a10870a  and  a10867a );
 a10874a <=( A232  and  (not A203) );
 a10878a <=( A268  and  A236 );
 a10879a <=( (not A233)  and  a10878a );
 a10880a <=( a10879a  and  a10874a );
 a10883a <=( A167  and  A168 );
 a10886a <=( A200  and  A199 );
 a10887a <=( a10886a  and  a10883a );
 a10890a <=( (not A202)  and  (not A201) );
 a10894a <=( A300  and  A299 );
 a10895a <=( A235  and  a10894a );
 a10896a <=( a10895a  and  a10890a );
 a10899a <=( A167  and  A168 );
 a10902a <=( A200  and  A199 );
 a10903a <=( a10902a  and  a10899a );
 a10906a <=( (not A202)  and  (not A201) );
 a10910a <=( A300  and  A298 );
 a10911a <=( A235  and  a10910a );
 a10912a <=( a10911a  and  a10906a );
 a10915a <=( A167  and  A168 );
 a10918a <=( A200  and  A199 );
 a10919a <=( a10918a  and  a10915a );
 a10922a <=( (not A202)  and  (not A201) );
 a10926a <=( A267  and  A265 );
 a10927a <=( A235  and  a10926a );
 a10928a <=( a10927a  and  a10922a );
 a10931a <=( A167  and  A168 );
 a10934a <=( A200  and  A199 );
 a10935a <=( a10934a  and  a10931a );
 a10938a <=( (not A202)  and  (not A201) );
 a10942a <=( A267  and  A266 );
 a10943a <=( A235  and  a10942a );
 a10944a <=( a10943a  and  a10938a );
 a10947a <=( A167  and  A168 );
 a10950a <=( A200  and  A199 );
 a10951a <=( a10950a  and  a10947a );
 a10954a <=( (not A202)  and  (not A201) );
 a10958a <=( A301  and  A234 );
 a10959a <=( A232  and  a10958a );
 a10960a <=( a10959a  and  a10954a );
 a10963a <=( A167  and  A168 );
 a10966a <=( A200  and  A199 );
 a10967a <=( a10966a  and  a10963a );
 a10970a <=( (not A202)  and  (not A201) );
 a10974a <=( A268  and  A234 );
 a10975a <=( A232  and  a10974a );
 a10976a <=( a10975a  and  a10970a );
 a10979a <=( A167  and  A168 );
 a10982a <=( A200  and  A199 );
 a10983a <=( a10982a  and  a10979a );
 a10986a <=( (not A202)  and  (not A201) );
 a10990a <=( A301  and  A234 );
 a10991a <=( A233  and  a10990a );
 a10992a <=( a10991a  and  a10986a );
 a10995a <=( A167  and  A168 );
 a10998a <=( A200  and  A199 );
 a10999a <=( a10998a  and  a10995a );
 a11002a <=( (not A202)  and  (not A201) );
 a11006a <=( A268  and  A234 );
 a11007a <=( A233  and  a11006a );
 a11008a <=( a11007a  and  a11002a );
 a11011a <=( A167  and  A168 );
 a11014a <=( (not A200)  and  (not A199) );
 a11015a <=( a11014a  and  a11011a );
 a11018a <=( A235  and  (not A202) );
 a11022a <=( A302  and  (not A299) );
 a11023a <=( A298  and  a11022a );
 a11024a <=( a11023a  and  a11018a );
 a11027a <=( A167  and  A168 );
 a11030a <=( (not A200)  and  (not A199) );
 a11031a <=( a11030a  and  a11027a );
 a11034a <=( A235  and  (not A202) );
 a11038a <=( A302  and  A299 );
 a11039a <=( (not A298)  and  a11038a );
 a11040a <=( a11039a  and  a11034a );
 a11043a <=( A167  and  A168 );
 a11046a <=( (not A200)  and  (not A199) );
 a11047a <=( a11046a  and  a11043a );
 a11050a <=( A235  and  (not A202) );
 a11054a <=( A269  and  A266 );
 a11055a <=( (not A265)  and  a11054a );
 a11056a <=( a11055a  and  a11050a );
 a11059a <=( A167  and  A168 );
 a11062a <=( (not A200)  and  (not A199) );
 a11063a <=( a11062a  and  a11059a );
 a11066a <=( A235  and  (not A202) );
 a11070a <=( A269  and  (not A266) );
 a11071a <=( A265  and  a11070a );
 a11072a <=( a11071a  and  a11066a );
 a11075a <=( A167  and  A168 );
 a11078a <=( (not A200)  and  (not A199) );
 a11079a <=( a11078a  and  a11075a );
 a11082a <=( A232  and  (not A202) );
 a11086a <=( A300  and  A299 );
 a11087a <=( A234  and  a11086a );
 a11088a <=( a11087a  and  a11082a );
 a11091a <=( A167  and  A168 );
 a11094a <=( (not A200)  and  (not A199) );
 a11095a <=( a11094a  and  a11091a );
 a11098a <=( A232  and  (not A202) );
 a11102a <=( A300  and  A298 );
 a11103a <=( A234  and  a11102a );
 a11104a <=( a11103a  and  a11098a );
 a11107a <=( A167  and  A168 );
 a11110a <=( (not A200)  and  (not A199) );
 a11111a <=( a11110a  and  a11107a );
 a11114a <=( A232  and  (not A202) );
 a11118a <=( A267  and  A265 );
 a11119a <=( A234  and  a11118a );
 a11120a <=( a11119a  and  a11114a );
 a11123a <=( A167  and  A168 );
 a11126a <=( (not A200)  and  (not A199) );
 a11127a <=( a11126a  and  a11123a );
 a11130a <=( A232  and  (not A202) );
 a11134a <=( A267  and  A266 );
 a11135a <=( A234  and  a11134a );
 a11136a <=( a11135a  and  a11130a );
 a11139a <=( A167  and  A168 );
 a11142a <=( (not A200)  and  (not A199) );
 a11143a <=( a11142a  and  a11139a );
 a11146a <=( A233  and  (not A202) );
 a11150a <=( A300  and  A299 );
 a11151a <=( A234  and  a11150a );
 a11152a <=( a11151a  and  a11146a );
 a11155a <=( A167  and  A168 );
 a11158a <=( (not A200)  and  (not A199) );
 a11159a <=( a11158a  and  a11155a );
 a11162a <=( A233  and  (not A202) );
 a11166a <=( A300  and  A298 );
 a11167a <=( A234  and  a11166a );
 a11168a <=( a11167a  and  a11162a );
 a11171a <=( A167  and  A168 );
 a11174a <=( (not A200)  and  (not A199) );
 a11175a <=( a11174a  and  a11171a );
 a11178a <=( A233  and  (not A202) );
 a11182a <=( A267  and  A265 );
 a11183a <=( A234  and  a11182a );
 a11184a <=( a11183a  and  a11178a );
 a11187a <=( A167  and  A168 );
 a11190a <=( (not A200)  and  (not A199) );
 a11191a <=( a11190a  and  a11187a );
 a11194a <=( A233  and  (not A202) );
 a11198a <=( A267  and  A266 );
 a11199a <=( A234  and  a11198a );
 a11200a <=( a11199a  and  a11194a );
 a11203a <=( A167  and  A168 );
 a11206a <=( (not A200)  and  (not A199) );
 a11207a <=( a11206a  and  a11203a );
 a11210a <=( (not A232)  and  (not A202) );
 a11214a <=( A301  and  A236 );
 a11215a <=( A233  and  a11214a );
 a11216a <=( a11215a  and  a11210a );
 a11219a <=( A167  and  A168 );
 a11222a <=( (not A200)  and  (not A199) );
 a11223a <=( a11222a  and  a11219a );
 a11226a <=( (not A232)  and  (not A202) );
 a11230a <=( A268  and  A236 );
 a11231a <=( A233  and  a11230a );
 a11232a <=( a11231a  and  a11226a );
 a11235a <=( A167  and  A168 );
 a11238a <=( (not A200)  and  (not A199) );
 a11239a <=( a11238a  and  a11235a );
 a11242a <=( A232  and  (not A202) );
 a11246a <=( A301  and  A236 );
 a11247a <=( (not A233)  and  a11246a );
 a11248a <=( a11247a  and  a11242a );
 a11251a <=( A167  and  A168 );
 a11254a <=( (not A200)  and  (not A199) );
 a11255a <=( a11254a  and  a11251a );
 a11258a <=( A232  and  (not A202) );
 a11262a <=( A268  and  A236 );
 a11263a <=( (not A233)  and  a11262a );
 a11264a <=( a11263a  and  a11258a );
 a11267a <=( A167  and  A170 );
 a11270a <=( (not A201)  and  (not A166) );
 a11271a <=( a11270a  and  a11267a );
 a11274a <=( (not A203)  and  (not A202) );
 a11278a <=( A300  and  A299 );
 a11279a <=( A235  and  a11278a );
 a11280a <=( a11279a  and  a11274a );
 a11283a <=( A167  and  A170 );
 a11286a <=( (not A201)  and  (not A166) );
 a11287a <=( a11286a  and  a11283a );
 a11290a <=( (not A203)  and  (not A202) );
 a11294a <=( A300  and  A298 );
 a11295a <=( A235  and  a11294a );
 a11296a <=( a11295a  and  a11290a );
 a11299a <=( A167  and  A170 );
 a11302a <=( (not A201)  and  (not A166) );
 a11303a <=( a11302a  and  a11299a );
 a11306a <=( (not A203)  and  (not A202) );
 a11310a <=( A267  and  A265 );
 a11311a <=( A235  and  a11310a );
 a11312a <=( a11311a  and  a11306a );
 a11315a <=( A167  and  A170 );
 a11318a <=( (not A201)  and  (not A166) );
 a11319a <=( a11318a  and  a11315a );
 a11322a <=( (not A203)  and  (not A202) );
 a11326a <=( A267  and  A266 );
 a11327a <=( A235  and  a11326a );
 a11328a <=( a11327a  and  a11322a );
 a11331a <=( A167  and  A170 );
 a11334a <=( (not A201)  and  (not A166) );
 a11335a <=( a11334a  and  a11331a );
 a11338a <=( (not A203)  and  (not A202) );
 a11342a <=( A301  and  A234 );
 a11343a <=( A232  and  a11342a );
 a11344a <=( a11343a  and  a11338a );
 a11347a <=( A167  and  A170 );
 a11350a <=( (not A201)  and  (not A166) );
 a11351a <=( a11350a  and  a11347a );
 a11354a <=( (not A203)  and  (not A202) );
 a11358a <=( A268  and  A234 );
 a11359a <=( A232  and  a11358a );
 a11360a <=( a11359a  and  a11354a );
 a11363a <=( A167  and  A170 );
 a11366a <=( (not A201)  and  (not A166) );
 a11367a <=( a11366a  and  a11363a );
 a11370a <=( (not A203)  and  (not A202) );
 a11374a <=( A301  and  A234 );
 a11375a <=( A233  and  a11374a );
 a11376a <=( a11375a  and  a11370a );
 a11379a <=( A167  and  A170 );
 a11382a <=( (not A201)  and  (not A166) );
 a11383a <=( a11382a  and  a11379a );
 a11386a <=( (not A203)  and  (not A202) );
 a11390a <=( A268  and  A234 );
 a11391a <=( A233  and  a11390a );
 a11392a <=( a11391a  and  a11386a );
 a11395a <=( A167  and  A170 );
 a11398a <=( A199  and  (not A166) );
 a11399a <=( a11398a  and  a11395a );
 a11402a <=( (not A201)  and  A200 );
 a11406a <=( A301  and  A235 );
 a11407a <=( (not A202)  and  a11406a );
 a11408a <=( a11407a  and  a11402a );
 a11411a <=( A167  and  A170 );
 a11414a <=( A199  and  (not A166) );
 a11415a <=( a11414a  and  a11411a );
 a11418a <=( (not A201)  and  A200 );
 a11422a <=( A268  and  A235 );
 a11423a <=( (not A202)  and  a11422a );
 a11424a <=( a11423a  and  a11418a );
 a11427a <=( A167  and  A170 );
 a11430a <=( (not A199)  and  (not A166) );
 a11431a <=( a11430a  and  a11427a );
 a11434a <=( (not A202)  and  (not A200) );
 a11438a <=( A300  and  A299 );
 a11439a <=( A235  and  a11438a );
 a11440a <=( a11439a  and  a11434a );
 a11443a <=( A167  and  A170 );
 a11446a <=( (not A199)  and  (not A166) );
 a11447a <=( a11446a  and  a11443a );
 a11450a <=( (not A202)  and  (not A200) );
 a11454a <=( A300  and  A298 );
 a11455a <=( A235  and  a11454a );
 a11456a <=( a11455a  and  a11450a );
 a11459a <=( A167  and  A170 );
 a11462a <=( (not A199)  and  (not A166) );
 a11463a <=( a11462a  and  a11459a );
 a11466a <=( (not A202)  and  (not A200) );
 a11470a <=( A267  and  A265 );
 a11471a <=( A235  and  a11470a );
 a11472a <=( a11471a  and  a11466a );
 a11475a <=( A167  and  A170 );
 a11478a <=( (not A199)  and  (not A166) );
 a11479a <=( a11478a  and  a11475a );
 a11482a <=( (not A202)  and  (not A200) );
 a11486a <=( A267  and  A266 );
 a11487a <=( A235  and  a11486a );
 a11488a <=( a11487a  and  a11482a );
 a11491a <=( A167  and  A170 );
 a11494a <=( (not A199)  and  (not A166) );
 a11495a <=( a11494a  and  a11491a );
 a11498a <=( (not A202)  and  (not A200) );
 a11502a <=( A301  and  A234 );
 a11503a <=( A232  and  a11502a );
 a11504a <=( a11503a  and  a11498a );
 a11507a <=( A167  and  A170 );
 a11510a <=( (not A199)  and  (not A166) );
 a11511a <=( a11510a  and  a11507a );
 a11514a <=( (not A202)  and  (not A200) );
 a11518a <=( A268  and  A234 );
 a11519a <=( A232  and  a11518a );
 a11520a <=( a11519a  and  a11514a );
 a11523a <=( A167  and  A170 );
 a11526a <=( (not A199)  and  (not A166) );
 a11527a <=( a11526a  and  a11523a );
 a11530a <=( (not A202)  and  (not A200) );
 a11534a <=( A301  and  A234 );
 a11535a <=( A233  and  a11534a );
 a11536a <=( a11535a  and  a11530a );
 a11539a <=( A167  and  A170 );
 a11542a <=( (not A199)  and  (not A166) );
 a11543a <=( a11542a  and  a11539a );
 a11546a <=( (not A202)  and  (not A200) );
 a11550a <=( A268  and  A234 );
 a11551a <=( A233  and  a11550a );
 a11552a <=( a11551a  and  a11546a );
 a11555a <=( (not A167)  and  A170 );
 a11558a <=( (not A201)  and  A166 );
 a11559a <=( a11558a  and  a11555a );
 a11562a <=( (not A203)  and  (not A202) );
 a11566a <=( A300  and  A299 );
 a11567a <=( A235  and  a11566a );
 a11568a <=( a11567a  and  a11562a );
 a11571a <=( (not A167)  and  A170 );
 a11574a <=( (not A201)  and  A166 );
 a11575a <=( a11574a  and  a11571a );
 a11578a <=( (not A203)  and  (not A202) );
 a11582a <=( A300  and  A298 );
 a11583a <=( A235  and  a11582a );
 a11584a <=( a11583a  and  a11578a );
 a11587a <=( (not A167)  and  A170 );
 a11590a <=( (not A201)  and  A166 );
 a11591a <=( a11590a  and  a11587a );
 a11594a <=( (not A203)  and  (not A202) );
 a11598a <=( A267  and  A265 );
 a11599a <=( A235  and  a11598a );
 a11600a <=( a11599a  and  a11594a );
 a11603a <=( (not A167)  and  A170 );
 a11606a <=( (not A201)  and  A166 );
 a11607a <=( a11606a  and  a11603a );
 a11610a <=( (not A203)  and  (not A202) );
 a11614a <=( A267  and  A266 );
 a11615a <=( A235  and  a11614a );
 a11616a <=( a11615a  and  a11610a );
 a11619a <=( (not A167)  and  A170 );
 a11622a <=( (not A201)  and  A166 );
 a11623a <=( a11622a  and  a11619a );
 a11626a <=( (not A203)  and  (not A202) );
 a11630a <=( A301  and  A234 );
 a11631a <=( A232  and  a11630a );
 a11632a <=( a11631a  and  a11626a );
 a11635a <=( (not A167)  and  A170 );
 a11638a <=( (not A201)  and  A166 );
 a11639a <=( a11638a  and  a11635a );
 a11642a <=( (not A203)  and  (not A202) );
 a11646a <=( A268  and  A234 );
 a11647a <=( A232  and  a11646a );
 a11648a <=( a11647a  and  a11642a );
 a11651a <=( (not A167)  and  A170 );
 a11654a <=( (not A201)  and  A166 );
 a11655a <=( a11654a  and  a11651a );
 a11658a <=( (not A203)  and  (not A202) );
 a11662a <=( A301  and  A234 );
 a11663a <=( A233  and  a11662a );
 a11664a <=( a11663a  and  a11658a );
 a11667a <=( (not A167)  and  A170 );
 a11670a <=( (not A201)  and  A166 );
 a11671a <=( a11670a  and  a11667a );
 a11674a <=( (not A203)  and  (not A202) );
 a11678a <=( A268  and  A234 );
 a11679a <=( A233  and  a11678a );
 a11680a <=( a11679a  and  a11674a );
 a11683a <=( (not A167)  and  A170 );
 a11686a <=( A199  and  A166 );
 a11687a <=( a11686a  and  a11683a );
 a11690a <=( (not A201)  and  A200 );
 a11694a <=( A301  and  A235 );
 a11695a <=( (not A202)  and  a11694a );
 a11696a <=( a11695a  and  a11690a );
 a11699a <=( (not A167)  and  A170 );
 a11702a <=( A199  and  A166 );
 a11703a <=( a11702a  and  a11699a );
 a11706a <=( (not A201)  and  A200 );
 a11710a <=( A268  and  A235 );
 a11711a <=( (not A202)  and  a11710a );
 a11712a <=( a11711a  and  a11706a );
 a11715a <=( (not A167)  and  A170 );
 a11718a <=( (not A199)  and  A166 );
 a11719a <=( a11718a  and  a11715a );
 a11722a <=( (not A202)  and  (not A200) );
 a11726a <=( A300  and  A299 );
 a11727a <=( A235  and  a11726a );
 a11728a <=( a11727a  and  a11722a );
 a11731a <=( (not A167)  and  A170 );
 a11734a <=( (not A199)  and  A166 );
 a11735a <=( a11734a  and  a11731a );
 a11738a <=( (not A202)  and  (not A200) );
 a11742a <=( A300  and  A298 );
 a11743a <=( A235  and  a11742a );
 a11744a <=( a11743a  and  a11738a );
 a11747a <=( (not A167)  and  A170 );
 a11750a <=( (not A199)  and  A166 );
 a11751a <=( a11750a  and  a11747a );
 a11754a <=( (not A202)  and  (not A200) );
 a11758a <=( A267  and  A265 );
 a11759a <=( A235  and  a11758a );
 a11760a <=( a11759a  and  a11754a );
 a11763a <=( (not A167)  and  A170 );
 a11766a <=( (not A199)  and  A166 );
 a11767a <=( a11766a  and  a11763a );
 a11770a <=( (not A202)  and  (not A200) );
 a11774a <=( A267  and  A266 );
 a11775a <=( A235  and  a11774a );
 a11776a <=( a11775a  and  a11770a );
 a11779a <=( (not A167)  and  A170 );
 a11782a <=( (not A199)  and  A166 );
 a11783a <=( a11782a  and  a11779a );
 a11786a <=( (not A202)  and  (not A200) );
 a11790a <=( A301  and  A234 );
 a11791a <=( A232  and  a11790a );
 a11792a <=( a11791a  and  a11786a );
 a11795a <=( (not A167)  and  A170 );
 a11798a <=( (not A199)  and  A166 );
 a11799a <=( a11798a  and  a11795a );
 a11802a <=( (not A202)  and  (not A200) );
 a11806a <=( A268  and  A234 );
 a11807a <=( A232  and  a11806a );
 a11808a <=( a11807a  and  a11802a );
 a11811a <=( (not A167)  and  A170 );
 a11814a <=( (not A199)  and  A166 );
 a11815a <=( a11814a  and  a11811a );
 a11818a <=( (not A202)  and  (not A200) );
 a11822a <=( A301  and  A234 );
 a11823a <=( A233  and  a11822a );
 a11824a <=( a11823a  and  a11818a );
 a11827a <=( (not A167)  and  A170 );
 a11830a <=( (not A199)  and  A166 );
 a11831a <=( a11830a  and  a11827a );
 a11834a <=( (not A202)  and  (not A200) );
 a11838a <=( A268  and  A234 );
 a11839a <=( A233  and  a11838a );
 a11840a <=( a11839a  and  a11834a );
 a11843a <=( (not A201)  and  A169 );
 a11846a <=( (not A203)  and  (not A202) );
 a11847a <=( a11846a  and  a11843a );
 a11850a <=( A234  and  A232 );
 a11854a <=( A302  and  (not A299) );
 a11855a <=( A298  and  a11854a );
 a11856a <=( a11855a  and  a11850a );
 a11859a <=( (not A201)  and  A169 );
 a11862a <=( (not A203)  and  (not A202) );
 a11863a <=( a11862a  and  a11859a );
 a11866a <=( A234  and  A232 );
 a11870a <=( A302  and  A299 );
 a11871a <=( (not A298)  and  a11870a );
 a11872a <=( a11871a  and  a11866a );
 a11875a <=( (not A201)  and  A169 );
 a11878a <=( (not A203)  and  (not A202) );
 a11879a <=( a11878a  and  a11875a );
 a11882a <=( A234  and  A232 );
 a11886a <=( A269  and  A266 );
 a11887a <=( (not A265)  and  a11886a );
 a11888a <=( a11887a  and  a11882a );
 a11891a <=( (not A201)  and  A169 );
 a11894a <=( (not A203)  and  (not A202) );
 a11895a <=( a11894a  and  a11891a );
 a11898a <=( A234  and  A232 );
 a11902a <=( A269  and  (not A266) );
 a11903a <=( A265  and  a11902a );
 a11904a <=( a11903a  and  a11898a );
 a11907a <=( (not A201)  and  A169 );
 a11910a <=( (not A203)  and  (not A202) );
 a11911a <=( a11910a  and  a11907a );
 a11914a <=( A234  and  A233 );
 a11918a <=( A302  and  (not A299) );
 a11919a <=( A298  and  a11918a );
 a11920a <=( a11919a  and  a11914a );
 a11923a <=( (not A201)  and  A169 );
 a11926a <=( (not A203)  and  (not A202) );
 a11927a <=( a11926a  and  a11923a );
 a11930a <=( A234  and  A233 );
 a11934a <=( A302  and  A299 );
 a11935a <=( (not A298)  and  a11934a );
 a11936a <=( a11935a  and  a11930a );
 a11939a <=( (not A201)  and  A169 );
 a11942a <=( (not A203)  and  (not A202) );
 a11943a <=( a11942a  and  a11939a );
 a11946a <=( A234  and  A233 );
 a11950a <=( A269  and  A266 );
 a11951a <=( (not A265)  and  a11950a );
 a11952a <=( a11951a  and  a11946a );
 a11955a <=( (not A201)  and  A169 );
 a11958a <=( (not A203)  and  (not A202) );
 a11959a <=( a11958a  and  a11955a );
 a11962a <=( A234  and  A233 );
 a11966a <=( A269  and  (not A266) );
 a11967a <=( A265  and  a11966a );
 a11968a <=( a11967a  and  a11962a );
 a11971a <=( (not A201)  and  A169 );
 a11974a <=( (not A203)  and  (not A202) );
 a11975a <=( a11974a  and  a11971a );
 a11978a <=( A233  and  (not A232) );
 a11982a <=( A300  and  A299 );
 a11983a <=( A236  and  a11982a );
 a11984a <=( a11983a  and  a11978a );
 a11987a <=( (not A201)  and  A169 );
 a11990a <=( (not A203)  and  (not A202) );
 a11991a <=( a11990a  and  a11987a );
 a11994a <=( A233  and  (not A232) );
 a11998a <=( A300  and  A298 );
 a11999a <=( A236  and  a11998a );
 a12000a <=( a11999a  and  a11994a );
 a12003a <=( (not A201)  and  A169 );
 a12006a <=( (not A203)  and  (not A202) );
 a12007a <=( a12006a  and  a12003a );
 a12010a <=( A233  and  (not A232) );
 a12014a <=( A267  and  A265 );
 a12015a <=( A236  and  a12014a );
 a12016a <=( a12015a  and  a12010a );
 a12019a <=( (not A201)  and  A169 );
 a12022a <=( (not A203)  and  (not A202) );
 a12023a <=( a12022a  and  a12019a );
 a12026a <=( A233  and  (not A232) );
 a12030a <=( A267  and  A266 );
 a12031a <=( A236  and  a12030a );
 a12032a <=( a12031a  and  a12026a );
 a12035a <=( (not A201)  and  A169 );
 a12038a <=( (not A203)  and  (not A202) );
 a12039a <=( a12038a  and  a12035a );
 a12042a <=( (not A233)  and  A232 );
 a12046a <=( A300  and  A299 );
 a12047a <=( A236  and  a12046a );
 a12048a <=( a12047a  and  a12042a );
 a12051a <=( (not A201)  and  A169 );
 a12054a <=( (not A203)  and  (not A202) );
 a12055a <=( a12054a  and  a12051a );
 a12058a <=( (not A233)  and  A232 );
 a12062a <=( A300  and  A298 );
 a12063a <=( A236  and  a12062a );
 a12064a <=( a12063a  and  a12058a );
 a12067a <=( (not A201)  and  A169 );
 a12070a <=( (not A203)  and  (not A202) );
 a12071a <=( a12070a  and  a12067a );
 a12074a <=( (not A233)  and  A232 );
 a12078a <=( A267  and  A265 );
 a12079a <=( A236  and  a12078a );
 a12080a <=( a12079a  and  a12074a );
 a12083a <=( (not A201)  and  A169 );
 a12086a <=( (not A203)  and  (not A202) );
 a12087a <=( a12086a  and  a12083a );
 a12090a <=( (not A233)  and  A232 );
 a12094a <=( A267  and  A266 );
 a12095a <=( A236  and  a12094a );
 a12096a <=( a12095a  and  a12090a );
 a12099a <=( A199  and  A169 );
 a12102a <=( (not A201)  and  A200 );
 a12103a <=( a12102a  and  a12099a );
 a12106a <=( A235  and  (not A202) );
 a12110a <=( A302  and  (not A299) );
 a12111a <=( A298  and  a12110a );
 a12112a <=( a12111a  and  a12106a );
 a12115a <=( A199  and  A169 );
 a12118a <=( (not A201)  and  A200 );
 a12119a <=( a12118a  and  a12115a );
 a12122a <=( A235  and  (not A202) );
 a12126a <=( A302  and  A299 );
 a12127a <=( (not A298)  and  a12126a );
 a12128a <=( a12127a  and  a12122a );
 a12131a <=( A199  and  A169 );
 a12134a <=( (not A201)  and  A200 );
 a12135a <=( a12134a  and  a12131a );
 a12138a <=( A235  and  (not A202) );
 a12142a <=( A269  and  A266 );
 a12143a <=( (not A265)  and  a12142a );
 a12144a <=( a12143a  and  a12138a );
 a12147a <=( A199  and  A169 );
 a12150a <=( (not A201)  and  A200 );
 a12151a <=( a12150a  and  a12147a );
 a12154a <=( A235  and  (not A202) );
 a12158a <=( A269  and  (not A266) );
 a12159a <=( A265  and  a12158a );
 a12160a <=( a12159a  and  a12154a );
 a12163a <=( A199  and  A169 );
 a12166a <=( (not A201)  and  A200 );
 a12167a <=( a12166a  and  a12163a );
 a12170a <=( A232  and  (not A202) );
 a12174a <=( A300  and  A299 );
 a12175a <=( A234  and  a12174a );
 a12176a <=( a12175a  and  a12170a );
 a12179a <=( A199  and  A169 );
 a12182a <=( (not A201)  and  A200 );
 a12183a <=( a12182a  and  a12179a );
 a12186a <=( A232  and  (not A202) );
 a12190a <=( A300  and  A298 );
 a12191a <=( A234  and  a12190a );
 a12192a <=( a12191a  and  a12186a );
 a12195a <=( A199  and  A169 );
 a12198a <=( (not A201)  and  A200 );
 a12199a <=( a12198a  and  a12195a );
 a12202a <=( A232  and  (not A202) );
 a12206a <=( A267  and  A265 );
 a12207a <=( A234  and  a12206a );
 a12208a <=( a12207a  and  a12202a );
 a12211a <=( A199  and  A169 );
 a12214a <=( (not A201)  and  A200 );
 a12215a <=( a12214a  and  a12211a );
 a12218a <=( A232  and  (not A202) );
 a12222a <=( A267  and  A266 );
 a12223a <=( A234  and  a12222a );
 a12224a <=( a12223a  and  a12218a );
 a12227a <=( A199  and  A169 );
 a12230a <=( (not A201)  and  A200 );
 a12231a <=( a12230a  and  a12227a );
 a12234a <=( A233  and  (not A202) );
 a12238a <=( A300  and  A299 );
 a12239a <=( A234  and  a12238a );
 a12240a <=( a12239a  and  a12234a );
 a12243a <=( A199  and  A169 );
 a12246a <=( (not A201)  and  A200 );
 a12247a <=( a12246a  and  a12243a );
 a12250a <=( A233  and  (not A202) );
 a12254a <=( A300  and  A298 );
 a12255a <=( A234  and  a12254a );
 a12256a <=( a12255a  and  a12250a );
 a12259a <=( A199  and  A169 );
 a12262a <=( (not A201)  and  A200 );
 a12263a <=( a12262a  and  a12259a );
 a12266a <=( A233  and  (not A202) );
 a12270a <=( A267  and  A265 );
 a12271a <=( A234  and  a12270a );
 a12272a <=( a12271a  and  a12266a );
 a12275a <=( A199  and  A169 );
 a12278a <=( (not A201)  and  A200 );
 a12279a <=( a12278a  and  a12275a );
 a12282a <=( A233  and  (not A202) );
 a12286a <=( A267  and  A266 );
 a12287a <=( A234  and  a12286a );
 a12288a <=( a12287a  and  a12282a );
 a12291a <=( A199  and  A169 );
 a12294a <=( (not A201)  and  A200 );
 a12295a <=( a12294a  and  a12291a );
 a12298a <=( (not A232)  and  (not A202) );
 a12302a <=( A301  and  A236 );
 a12303a <=( A233  and  a12302a );
 a12304a <=( a12303a  and  a12298a );
 a12307a <=( A199  and  A169 );
 a12310a <=( (not A201)  and  A200 );
 a12311a <=( a12310a  and  a12307a );
 a12314a <=( (not A232)  and  (not A202) );
 a12318a <=( A268  and  A236 );
 a12319a <=( A233  and  a12318a );
 a12320a <=( a12319a  and  a12314a );
 a12323a <=( A199  and  A169 );
 a12326a <=( (not A201)  and  A200 );
 a12327a <=( a12326a  and  a12323a );
 a12330a <=( A232  and  (not A202) );
 a12334a <=( A301  and  A236 );
 a12335a <=( (not A233)  and  a12334a );
 a12336a <=( a12335a  and  a12330a );
 a12339a <=( A199  and  A169 );
 a12342a <=( (not A201)  and  A200 );
 a12343a <=( a12342a  and  a12339a );
 a12346a <=( A232  and  (not A202) );
 a12350a <=( A268  and  A236 );
 a12351a <=( (not A233)  and  a12350a );
 a12352a <=( a12351a  and  a12346a );
 a12355a <=( (not A199)  and  A169 );
 a12358a <=( (not A202)  and  (not A200) );
 a12359a <=( a12358a  and  a12355a );
 a12362a <=( A234  and  A232 );
 a12366a <=( A302  and  (not A299) );
 a12367a <=( A298  and  a12366a );
 a12368a <=( a12367a  and  a12362a );
 a12371a <=( (not A199)  and  A169 );
 a12374a <=( (not A202)  and  (not A200) );
 a12375a <=( a12374a  and  a12371a );
 a12378a <=( A234  and  A232 );
 a12382a <=( A302  and  A299 );
 a12383a <=( (not A298)  and  a12382a );
 a12384a <=( a12383a  and  a12378a );
 a12387a <=( (not A199)  and  A169 );
 a12390a <=( (not A202)  and  (not A200) );
 a12391a <=( a12390a  and  a12387a );
 a12394a <=( A234  and  A232 );
 a12398a <=( A269  and  A266 );
 a12399a <=( (not A265)  and  a12398a );
 a12400a <=( a12399a  and  a12394a );
 a12403a <=( (not A199)  and  A169 );
 a12406a <=( (not A202)  and  (not A200) );
 a12407a <=( a12406a  and  a12403a );
 a12410a <=( A234  and  A232 );
 a12414a <=( A269  and  (not A266) );
 a12415a <=( A265  and  a12414a );
 a12416a <=( a12415a  and  a12410a );
 a12419a <=( (not A199)  and  A169 );
 a12422a <=( (not A202)  and  (not A200) );
 a12423a <=( a12422a  and  a12419a );
 a12426a <=( A234  and  A233 );
 a12430a <=( A302  and  (not A299) );
 a12431a <=( A298  and  a12430a );
 a12432a <=( a12431a  and  a12426a );
 a12435a <=( (not A199)  and  A169 );
 a12438a <=( (not A202)  and  (not A200) );
 a12439a <=( a12438a  and  a12435a );
 a12442a <=( A234  and  A233 );
 a12446a <=( A302  and  A299 );
 a12447a <=( (not A298)  and  a12446a );
 a12448a <=( a12447a  and  a12442a );
 a12451a <=( (not A199)  and  A169 );
 a12454a <=( (not A202)  and  (not A200) );
 a12455a <=( a12454a  and  a12451a );
 a12458a <=( A234  and  A233 );
 a12462a <=( A269  and  A266 );
 a12463a <=( (not A265)  and  a12462a );
 a12464a <=( a12463a  and  a12458a );
 a12467a <=( (not A199)  and  A169 );
 a12470a <=( (not A202)  and  (not A200) );
 a12471a <=( a12470a  and  a12467a );
 a12474a <=( A234  and  A233 );
 a12478a <=( A269  and  (not A266) );
 a12479a <=( A265  and  a12478a );
 a12480a <=( a12479a  and  a12474a );
 a12483a <=( (not A199)  and  A169 );
 a12486a <=( (not A202)  and  (not A200) );
 a12487a <=( a12486a  and  a12483a );
 a12490a <=( A233  and  (not A232) );
 a12494a <=( A300  and  A299 );
 a12495a <=( A236  and  a12494a );
 a12496a <=( a12495a  and  a12490a );
 a12499a <=( (not A199)  and  A169 );
 a12502a <=( (not A202)  and  (not A200) );
 a12503a <=( a12502a  and  a12499a );
 a12506a <=( A233  and  (not A232) );
 a12510a <=( A300  and  A298 );
 a12511a <=( A236  and  a12510a );
 a12512a <=( a12511a  and  a12506a );
 a12515a <=( (not A199)  and  A169 );
 a12518a <=( (not A202)  and  (not A200) );
 a12519a <=( a12518a  and  a12515a );
 a12522a <=( A233  and  (not A232) );
 a12526a <=( A267  and  A265 );
 a12527a <=( A236  and  a12526a );
 a12528a <=( a12527a  and  a12522a );
 a12531a <=( (not A199)  and  A169 );
 a12534a <=( (not A202)  and  (not A200) );
 a12535a <=( a12534a  and  a12531a );
 a12538a <=( A233  and  (not A232) );
 a12542a <=( A267  and  A266 );
 a12543a <=( A236  and  a12542a );
 a12544a <=( a12543a  and  a12538a );
 a12547a <=( (not A199)  and  A169 );
 a12550a <=( (not A202)  and  (not A200) );
 a12551a <=( a12550a  and  a12547a );
 a12554a <=( (not A233)  and  A232 );
 a12558a <=( A300  and  A299 );
 a12559a <=( A236  and  a12558a );
 a12560a <=( a12559a  and  a12554a );
 a12563a <=( (not A199)  and  A169 );
 a12566a <=( (not A202)  and  (not A200) );
 a12567a <=( a12566a  and  a12563a );
 a12570a <=( (not A233)  and  A232 );
 a12574a <=( A300  and  A298 );
 a12575a <=( A236  and  a12574a );
 a12576a <=( a12575a  and  a12570a );
 a12579a <=( (not A199)  and  A169 );
 a12582a <=( (not A202)  and  (not A200) );
 a12583a <=( a12582a  and  a12579a );
 a12586a <=( (not A233)  and  A232 );
 a12590a <=( A267  and  A265 );
 a12591a <=( A236  and  a12590a );
 a12592a <=( a12591a  and  a12586a );
 a12595a <=( (not A199)  and  A169 );
 a12598a <=( (not A202)  and  (not A200) );
 a12599a <=( a12598a  and  a12595a );
 a12602a <=( (not A233)  and  A232 );
 a12606a <=( A267  and  A266 );
 a12607a <=( A236  and  a12606a );
 a12608a <=( a12607a  and  a12602a );
 a12611a <=( (not A167)  and  (not A169) );
 a12614a <=( A202  and  (not A166) );
 a12615a <=( a12614a  and  a12611a );
 a12618a <=( A234  and  A232 );
 a12622a <=( A302  and  (not A299) );
 a12623a <=( A298  and  a12622a );
 a12624a <=( a12623a  and  a12618a );
 a12627a <=( (not A167)  and  (not A169) );
 a12630a <=( A202  and  (not A166) );
 a12631a <=( a12630a  and  a12627a );
 a12634a <=( A234  and  A232 );
 a12638a <=( A302  and  A299 );
 a12639a <=( (not A298)  and  a12638a );
 a12640a <=( a12639a  and  a12634a );
 a12643a <=( (not A167)  and  (not A169) );
 a12646a <=( A202  and  (not A166) );
 a12647a <=( a12646a  and  a12643a );
 a12650a <=( A234  and  A232 );
 a12654a <=( A269  and  A266 );
 a12655a <=( (not A265)  and  a12654a );
 a12656a <=( a12655a  and  a12650a );
 a12659a <=( (not A167)  and  (not A169) );
 a12662a <=( A202  and  (not A166) );
 a12663a <=( a12662a  and  a12659a );
 a12666a <=( A234  and  A232 );
 a12670a <=( A269  and  (not A266) );
 a12671a <=( A265  and  a12670a );
 a12672a <=( a12671a  and  a12666a );
 a12675a <=( (not A167)  and  (not A169) );
 a12678a <=( A202  and  (not A166) );
 a12679a <=( a12678a  and  a12675a );
 a12682a <=( A234  and  A233 );
 a12686a <=( A302  and  (not A299) );
 a12687a <=( A298  and  a12686a );
 a12688a <=( a12687a  and  a12682a );
 a12691a <=( (not A167)  and  (not A169) );
 a12694a <=( A202  and  (not A166) );
 a12695a <=( a12694a  and  a12691a );
 a12698a <=( A234  and  A233 );
 a12702a <=( A302  and  A299 );
 a12703a <=( (not A298)  and  a12702a );
 a12704a <=( a12703a  and  a12698a );
 a12707a <=( (not A167)  and  (not A169) );
 a12710a <=( A202  and  (not A166) );
 a12711a <=( a12710a  and  a12707a );
 a12714a <=( A234  and  A233 );
 a12718a <=( A269  and  A266 );
 a12719a <=( (not A265)  and  a12718a );
 a12720a <=( a12719a  and  a12714a );
 a12723a <=( (not A167)  and  (not A169) );
 a12726a <=( A202  and  (not A166) );
 a12727a <=( a12726a  and  a12723a );
 a12730a <=( A234  and  A233 );
 a12734a <=( A269  and  (not A266) );
 a12735a <=( A265  and  a12734a );
 a12736a <=( a12735a  and  a12730a );
 a12739a <=( (not A167)  and  (not A169) );
 a12742a <=( A202  and  (not A166) );
 a12743a <=( a12742a  and  a12739a );
 a12746a <=( A233  and  (not A232) );
 a12750a <=( A300  and  A299 );
 a12751a <=( A236  and  a12750a );
 a12752a <=( a12751a  and  a12746a );
 a12755a <=( (not A167)  and  (not A169) );
 a12758a <=( A202  and  (not A166) );
 a12759a <=( a12758a  and  a12755a );
 a12762a <=( A233  and  (not A232) );
 a12766a <=( A300  and  A298 );
 a12767a <=( A236  and  a12766a );
 a12768a <=( a12767a  and  a12762a );
 a12771a <=( (not A167)  and  (not A169) );
 a12774a <=( A202  and  (not A166) );
 a12775a <=( a12774a  and  a12771a );
 a12778a <=( A233  and  (not A232) );
 a12782a <=( A267  and  A265 );
 a12783a <=( A236  and  a12782a );
 a12784a <=( a12783a  and  a12778a );
 a12787a <=( (not A167)  and  (not A169) );
 a12790a <=( A202  and  (not A166) );
 a12791a <=( a12790a  and  a12787a );
 a12794a <=( A233  and  (not A232) );
 a12798a <=( A267  and  A266 );
 a12799a <=( A236  and  a12798a );
 a12800a <=( a12799a  and  a12794a );
 a12803a <=( (not A167)  and  (not A169) );
 a12806a <=( A202  and  (not A166) );
 a12807a <=( a12806a  and  a12803a );
 a12810a <=( (not A233)  and  A232 );
 a12814a <=( A300  and  A299 );
 a12815a <=( A236  and  a12814a );
 a12816a <=( a12815a  and  a12810a );
 a12819a <=( (not A167)  and  (not A169) );
 a12822a <=( A202  and  (not A166) );
 a12823a <=( a12822a  and  a12819a );
 a12826a <=( (not A233)  and  A232 );
 a12830a <=( A300  and  A298 );
 a12831a <=( A236  and  a12830a );
 a12832a <=( a12831a  and  a12826a );
 a12835a <=( (not A167)  and  (not A169) );
 a12838a <=( A202  and  (not A166) );
 a12839a <=( a12838a  and  a12835a );
 a12842a <=( (not A233)  and  A232 );
 a12846a <=( A267  and  A265 );
 a12847a <=( A236  and  a12846a );
 a12848a <=( a12847a  and  a12842a );
 a12851a <=( (not A167)  and  (not A169) );
 a12854a <=( A202  and  (not A166) );
 a12855a <=( a12854a  and  a12851a );
 a12858a <=( (not A233)  and  A232 );
 a12862a <=( A267  and  A266 );
 a12863a <=( A236  and  a12862a );
 a12864a <=( a12863a  and  a12858a );
 a12867a <=( (not A167)  and  (not A169) );
 a12870a <=( A199  and  (not A166) );
 a12871a <=( a12870a  and  a12867a );
 a12874a <=( A235  and  A201 );
 a12878a <=( A302  and  (not A299) );
 a12879a <=( A298  and  a12878a );
 a12880a <=( a12879a  and  a12874a );
 a12883a <=( (not A167)  and  (not A169) );
 a12886a <=( A199  and  (not A166) );
 a12887a <=( a12886a  and  a12883a );
 a12890a <=( A235  and  A201 );
 a12894a <=( A302  and  A299 );
 a12895a <=( (not A298)  and  a12894a );
 a12896a <=( a12895a  and  a12890a );
 a12899a <=( (not A167)  and  (not A169) );
 a12902a <=( A199  and  (not A166) );
 a12903a <=( a12902a  and  a12899a );
 a12906a <=( A235  and  A201 );
 a12910a <=( A269  and  A266 );
 a12911a <=( (not A265)  and  a12910a );
 a12912a <=( a12911a  and  a12906a );
 a12915a <=( (not A167)  and  (not A169) );
 a12918a <=( A199  and  (not A166) );
 a12919a <=( a12918a  and  a12915a );
 a12922a <=( A235  and  A201 );
 a12926a <=( A269  and  (not A266) );
 a12927a <=( A265  and  a12926a );
 a12928a <=( a12927a  and  a12922a );
 a12931a <=( (not A167)  and  (not A169) );
 a12934a <=( A199  and  (not A166) );
 a12935a <=( a12934a  and  a12931a );
 a12938a <=( A232  and  A201 );
 a12942a <=( A300  and  A299 );
 a12943a <=( A234  and  a12942a );
 a12944a <=( a12943a  and  a12938a );
 a12947a <=( (not A167)  and  (not A169) );
 a12950a <=( A199  and  (not A166) );
 a12951a <=( a12950a  and  a12947a );
 a12954a <=( A232  and  A201 );
 a12958a <=( A300  and  A298 );
 a12959a <=( A234  and  a12958a );
 a12960a <=( a12959a  and  a12954a );
 a12963a <=( (not A167)  and  (not A169) );
 a12966a <=( A199  and  (not A166) );
 a12967a <=( a12966a  and  a12963a );
 a12970a <=( A232  and  A201 );
 a12974a <=( A267  and  A265 );
 a12975a <=( A234  and  a12974a );
 a12976a <=( a12975a  and  a12970a );
 a12979a <=( (not A167)  and  (not A169) );
 a12982a <=( A199  and  (not A166) );
 a12983a <=( a12982a  and  a12979a );
 a12986a <=( A232  and  A201 );
 a12990a <=( A267  and  A266 );
 a12991a <=( A234  and  a12990a );
 a12992a <=( a12991a  and  a12986a );
 a12995a <=( (not A167)  and  (not A169) );
 a12998a <=( A199  and  (not A166) );
 a12999a <=( a12998a  and  a12995a );
 a13002a <=( A233  and  A201 );
 a13006a <=( A300  and  A299 );
 a13007a <=( A234  and  a13006a );
 a13008a <=( a13007a  and  a13002a );
 a13011a <=( (not A167)  and  (not A169) );
 a13014a <=( A199  and  (not A166) );
 a13015a <=( a13014a  and  a13011a );
 a13018a <=( A233  and  A201 );
 a13022a <=( A300  and  A298 );
 a13023a <=( A234  and  a13022a );
 a13024a <=( a13023a  and  a13018a );
 a13027a <=( (not A167)  and  (not A169) );
 a13030a <=( A199  and  (not A166) );
 a13031a <=( a13030a  and  a13027a );
 a13034a <=( A233  and  A201 );
 a13038a <=( A267  and  A265 );
 a13039a <=( A234  and  a13038a );
 a13040a <=( a13039a  and  a13034a );
 a13043a <=( (not A167)  and  (not A169) );
 a13046a <=( A199  and  (not A166) );
 a13047a <=( a13046a  and  a13043a );
 a13050a <=( A233  and  A201 );
 a13054a <=( A267  and  A266 );
 a13055a <=( A234  and  a13054a );
 a13056a <=( a13055a  and  a13050a );
 a13059a <=( (not A167)  and  (not A169) );
 a13062a <=( A199  and  (not A166) );
 a13063a <=( a13062a  and  a13059a );
 a13066a <=( (not A232)  and  A201 );
 a13070a <=( A301  and  A236 );
 a13071a <=( A233  and  a13070a );
 a13072a <=( a13071a  and  a13066a );
 a13075a <=( (not A167)  and  (not A169) );
 a13078a <=( A199  and  (not A166) );
 a13079a <=( a13078a  and  a13075a );
 a13082a <=( (not A232)  and  A201 );
 a13086a <=( A268  and  A236 );
 a13087a <=( A233  and  a13086a );
 a13088a <=( a13087a  and  a13082a );
 a13091a <=( (not A167)  and  (not A169) );
 a13094a <=( A199  and  (not A166) );
 a13095a <=( a13094a  and  a13091a );
 a13098a <=( A232  and  A201 );
 a13102a <=( A301  and  A236 );
 a13103a <=( (not A233)  and  a13102a );
 a13104a <=( a13103a  and  a13098a );
 a13107a <=( (not A167)  and  (not A169) );
 a13110a <=( A199  and  (not A166) );
 a13111a <=( a13110a  and  a13107a );
 a13114a <=( A232  and  A201 );
 a13118a <=( A268  and  A236 );
 a13119a <=( (not A233)  and  a13118a );
 a13120a <=( a13119a  and  a13114a );
 a13123a <=( (not A167)  and  (not A169) );
 a13126a <=( A200  and  (not A166) );
 a13127a <=( a13126a  and  a13123a );
 a13130a <=( A235  and  A201 );
 a13134a <=( A302  and  (not A299) );
 a13135a <=( A298  and  a13134a );
 a13136a <=( a13135a  and  a13130a );
 a13139a <=( (not A167)  and  (not A169) );
 a13142a <=( A200  and  (not A166) );
 a13143a <=( a13142a  and  a13139a );
 a13146a <=( A235  and  A201 );
 a13150a <=( A302  and  A299 );
 a13151a <=( (not A298)  and  a13150a );
 a13152a <=( a13151a  and  a13146a );
 a13155a <=( (not A167)  and  (not A169) );
 a13158a <=( A200  and  (not A166) );
 a13159a <=( a13158a  and  a13155a );
 a13162a <=( A235  and  A201 );
 a13166a <=( A269  and  A266 );
 a13167a <=( (not A265)  and  a13166a );
 a13168a <=( a13167a  and  a13162a );
 a13171a <=( (not A167)  and  (not A169) );
 a13174a <=( A200  and  (not A166) );
 a13175a <=( a13174a  and  a13171a );
 a13178a <=( A235  and  A201 );
 a13182a <=( A269  and  (not A266) );
 a13183a <=( A265  and  a13182a );
 a13184a <=( a13183a  and  a13178a );
 a13187a <=( (not A167)  and  (not A169) );
 a13190a <=( A200  and  (not A166) );
 a13191a <=( a13190a  and  a13187a );
 a13194a <=( A232  and  A201 );
 a13198a <=( A300  and  A299 );
 a13199a <=( A234  and  a13198a );
 a13200a <=( a13199a  and  a13194a );
 a13203a <=( (not A167)  and  (not A169) );
 a13206a <=( A200  and  (not A166) );
 a13207a <=( a13206a  and  a13203a );
 a13210a <=( A232  and  A201 );
 a13214a <=( A300  and  A298 );
 a13215a <=( A234  and  a13214a );
 a13216a <=( a13215a  and  a13210a );
 a13219a <=( (not A167)  and  (not A169) );
 a13222a <=( A200  and  (not A166) );
 a13223a <=( a13222a  and  a13219a );
 a13226a <=( A232  and  A201 );
 a13230a <=( A267  and  A265 );
 a13231a <=( A234  and  a13230a );
 a13232a <=( a13231a  and  a13226a );
 a13235a <=( (not A167)  and  (not A169) );
 a13238a <=( A200  and  (not A166) );
 a13239a <=( a13238a  and  a13235a );
 a13242a <=( A232  and  A201 );
 a13246a <=( A267  and  A266 );
 a13247a <=( A234  and  a13246a );
 a13248a <=( a13247a  and  a13242a );
 a13251a <=( (not A167)  and  (not A169) );
 a13254a <=( A200  and  (not A166) );
 a13255a <=( a13254a  and  a13251a );
 a13258a <=( A233  and  A201 );
 a13262a <=( A300  and  A299 );
 a13263a <=( A234  and  a13262a );
 a13264a <=( a13263a  and  a13258a );
 a13267a <=( (not A167)  and  (not A169) );
 a13270a <=( A200  and  (not A166) );
 a13271a <=( a13270a  and  a13267a );
 a13274a <=( A233  and  A201 );
 a13278a <=( A300  and  A298 );
 a13279a <=( A234  and  a13278a );
 a13280a <=( a13279a  and  a13274a );
 a13283a <=( (not A167)  and  (not A169) );
 a13286a <=( A200  and  (not A166) );
 a13287a <=( a13286a  and  a13283a );
 a13290a <=( A233  and  A201 );
 a13294a <=( A267  and  A265 );
 a13295a <=( A234  and  a13294a );
 a13296a <=( a13295a  and  a13290a );
 a13299a <=( (not A167)  and  (not A169) );
 a13302a <=( A200  and  (not A166) );
 a13303a <=( a13302a  and  a13299a );
 a13306a <=( A233  and  A201 );
 a13310a <=( A267  and  A266 );
 a13311a <=( A234  and  a13310a );
 a13312a <=( a13311a  and  a13306a );
 a13315a <=( (not A167)  and  (not A169) );
 a13318a <=( A200  and  (not A166) );
 a13319a <=( a13318a  and  a13315a );
 a13322a <=( (not A232)  and  A201 );
 a13326a <=( A301  and  A236 );
 a13327a <=( A233  and  a13326a );
 a13328a <=( a13327a  and  a13322a );
 a13331a <=( (not A167)  and  (not A169) );
 a13334a <=( A200  and  (not A166) );
 a13335a <=( a13334a  and  a13331a );
 a13338a <=( (not A232)  and  A201 );
 a13342a <=( A268  and  A236 );
 a13343a <=( A233  and  a13342a );
 a13344a <=( a13343a  and  a13338a );
 a13347a <=( (not A167)  and  (not A169) );
 a13350a <=( A200  and  (not A166) );
 a13351a <=( a13350a  and  a13347a );
 a13354a <=( A232  and  A201 );
 a13358a <=( A301  and  A236 );
 a13359a <=( (not A233)  and  a13358a );
 a13360a <=( a13359a  and  a13354a );
 a13363a <=( (not A167)  and  (not A169) );
 a13366a <=( A200  and  (not A166) );
 a13367a <=( a13366a  and  a13363a );
 a13370a <=( A232  and  A201 );
 a13374a <=( A268  and  A236 );
 a13375a <=( (not A233)  and  a13374a );
 a13376a <=( a13375a  and  a13370a );
 a13379a <=( (not A167)  and  (not A169) );
 a13382a <=( (not A199)  and  (not A166) );
 a13383a <=( a13382a  and  a13379a );
 a13386a <=( A203  and  A200 );
 a13390a <=( A300  and  A299 );
 a13391a <=( A235  and  a13390a );
 a13392a <=( a13391a  and  a13386a );
 a13395a <=( (not A167)  and  (not A169) );
 a13398a <=( (not A199)  and  (not A166) );
 a13399a <=( a13398a  and  a13395a );
 a13402a <=( A203  and  A200 );
 a13406a <=( A300  and  A298 );
 a13407a <=( A235  and  a13406a );
 a13408a <=( a13407a  and  a13402a );
 a13411a <=( (not A167)  and  (not A169) );
 a13414a <=( (not A199)  and  (not A166) );
 a13415a <=( a13414a  and  a13411a );
 a13418a <=( A203  and  A200 );
 a13422a <=( A267  and  A265 );
 a13423a <=( A235  and  a13422a );
 a13424a <=( a13423a  and  a13418a );
 a13427a <=( (not A167)  and  (not A169) );
 a13430a <=( (not A199)  and  (not A166) );
 a13431a <=( a13430a  and  a13427a );
 a13434a <=( A203  and  A200 );
 a13438a <=( A267  and  A266 );
 a13439a <=( A235  and  a13438a );
 a13440a <=( a13439a  and  a13434a );
 a13443a <=( (not A167)  and  (not A169) );
 a13446a <=( (not A199)  and  (not A166) );
 a13447a <=( a13446a  and  a13443a );
 a13450a <=( A203  and  A200 );
 a13454a <=( A301  and  A234 );
 a13455a <=( A232  and  a13454a );
 a13456a <=( a13455a  and  a13450a );
 a13459a <=( (not A167)  and  (not A169) );
 a13462a <=( (not A199)  and  (not A166) );
 a13463a <=( a13462a  and  a13459a );
 a13466a <=( A203  and  A200 );
 a13470a <=( A268  and  A234 );
 a13471a <=( A232  and  a13470a );
 a13472a <=( a13471a  and  a13466a );
 a13475a <=( (not A167)  and  (not A169) );
 a13478a <=( (not A199)  and  (not A166) );
 a13479a <=( a13478a  and  a13475a );
 a13482a <=( A203  and  A200 );
 a13486a <=( A301  and  A234 );
 a13487a <=( A233  and  a13486a );
 a13488a <=( a13487a  and  a13482a );
 a13491a <=( (not A167)  and  (not A169) );
 a13494a <=( (not A199)  and  (not A166) );
 a13495a <=( a13494a  and  a13491a );
 a13498a <=( A203  and  A200 );
 a13502a <=( A268  and  A234 );
 a13503a <=( A233  and  a13502a );
 a13504a <=( a13503a  and  a13498a );
 a13507a <=( (not A167)  and  (not A169) );
 a13510a <=( A199  and  (not A166) );
 a13511a <=( a13510a  and  a13507a );
 a13514a <=( A203  and  (not A200) );
 a13518a <=( A300  and  A299 );
 a13519a <=( A235  and  a13518a );
 a13520a <=( a13519a  and  a13514a );
 a13523a <=( (not A167)  and  (not A169) );
 a13526a <=( A199  and  (not A166) );
 a13527a <=( a13526a  and  a13523a );
 a13530a <=( A203  and  (not A200) );
 a13534a <=( A300  and  A298 );
 a13535a <=( A235  and  a13534a );
 a13536a <=( a13535a  and  a13530a );
 a13539a <=( (not A167)  and  (not A169) );
 a13542a <=( A199  and  (not A166) );
 a13543a <=( a13542a  and  a13539a );
 a13546a <=( A203  and  (not A200) );
 a13550a <=( A267  and  A265 );
 a13551a <=( A235  and  a13550a );
 a13552a <=( a13551a  and  a13546a );
 a13555a <=( (not A167)  and  (not A169) );
 a13558a <=( A199  and  (not A166) );
 a13559a <=( a13558a  and  a13555a );
 a13562a <=( A203  and  (not A200) );
 a13566a <=( A267  and  A266 );
 a13567a <=( A235  and  a13566a );
 a13568a <=( a13567a  and  a13562a );
 a13571a <=( (not A167)  and  (not A169) );
 a13574a <=( A199  and  (not A166) );
 a13575a <=( a13574a  and  a13571a );
 a13578a <=( A203  and  (not A200) );
 a13582a <=( A301  and  A234 );
 a13583a <=( A232  and  a13582a );
 a13584a <=( a13583a  and  a13578a );
 a13587a <=( (not A167)  and  (not A169) );
 a13590a <=( A199  and  (not A166) );
 a13591a <=( a13590a  and  a13587a );
 a13594a <=( A203  and  (not A200) );
 a13598a <=( A268  and  A234 );
 a13599a <=( A232  and  a13598a );
 a13600a <=( a13599a  and  a13594a );
 a13603a <=( (not A167)  and  (not A169) );
 a13606a <=( A199  and  (not A166) );
 a13607a <=( a13606a  and  a13603a );
 a13610a <=( A203  and  (not A200) );
 a13614a <=( A301  and  A234 );
 a13615a <=( A233  and  a13614a );
 a13616a <=( a13615a  and  a13610a );
 a13619a <=( (not A167)  and  (not A169) );
 a13622a <=( A199  and  (not A166) );
 a13623a <=( a13622a  and  a13619a );
 a13626a <=( A203  and  (not A200) );
 a13630a <=( A268  and  A234 );
 a13631a <=( A233  and  a13630a );
 a13632a <=( a13631a  and  a13626a );
 a13635a <=( (not A168)  and  (not A169) );
 a13638a <=( A166  and  A167 );
 a13639a <=( a13638a  and  a13635a );
 a13642a <=( A235  and  A202 );
 a13646a <=( A302  and  (not A299) );
 a13647a <=( A298  and  a13646a );
 a13648a <=( a13647a  and  a13642a );
 a13651a <=( (not A168)  and  (not A169) );
 a13654a <=( A166  and  A167 );
 a13655a <=( a13654a  and  a13651a );
 a13658a <=( A235  and  A202 );
 a13662a <=( A302  and  A299 );
 a13663a <=( (not A298)  and  a13662a );
 a13664a <=( a13663a  and  a13658a );
 a13667a <=( (not A168)  and  (not A169) );
 a13670a <=( A166  and  A167 );
 a13671a <=( a13670a  and  a13667a );
 a13674a <=( A235  and  A202 );
 a13678a <=( A269  and  A266 );
 a13679a <=( (not A265)  and  a13678a );
 a13680a <=( a13679a  and  a13674a );
 a13683a <=( (not A168)  and  (not A169) );
 a13686a <=( A166  and  A167 );
 a13687a <=( a13686a  and  a13683a );
 a13690a <=( A235  and  A202 );
 a13694a <=( A269  and  (not A266) );
 a13695a <=( A265  and  a13694a );
 a13696a <=( a13695a  and  a13690a );
 a13699a <=( (not A168)  and  (not A169) );
 a13702a <=( A166  and  A167 );
 a13703a <=( a13702a  and  a13699a );
 a13706a <=( A232  and  A202 );
 a13710a <=( A300  and  A299 );
 a13711a <=( A234  and  a13710a );
 a13712a <=( a13711a  and  a13706a );
 a13715a <=( (not A168)  and  (not A169) );
 a13718a <=( A166  and  A167 );
 a13719a <=( a13718a  and  a13715a );
 a13722a <=( A232  and  A202 );
 a13726a <=( A300  and  A298 );
 a13727a <=( A234  and  a13726a );
 a13728a <=( a13727a  and  a13722a );
 a13731a <=( (not A168)  and  (not A169) );
 a13734a <=( A166  and  A167 );
 a13735a <=( a13734a  and  a13731a );
 a13738a <=( A232  and  A202 );
 a13742a <=( A267  and  A265 );
 a13743a <=( A234  and  a13742a );
 a13744a <=( a13743a  and  a13738a );
 a13747a <=( (not A168)  and  (not A169) );
 a13750a <=( A166  and  A167 );
 a13751a <=( a13750a  and  a13747a );
 a13754a <=( A232  and  A202 );
 a13758a <=( A267  and  A266 );
 a13759a <=( A234  and  a13758a );
 a13760a <=( a13759a  and  a13754a );
 a13763a <=( (not A168)  and  (not A169) );
 a13766a <=( A166  and  A167 );
 a13767a <=( a13766a  and  a13763a );
 a13770a <=( A233  and  A202 );
 a13774a <=( A300  and  A299 );
 a13775a <=( A234  and  a13774a );
 a13776a <=( a13775a  and  a13770a );
 a13779a <=( (not A168)  and  (not A169) );
 a13782a <=( A166  and  A167 );
 a13783a <=( a13782a  and  a13779a );
 a13786a <=( A233  and  A202 );
 a13790a <=( A300  and  A298 );
 a13791a <=( A234  and  a13790a );
 a13792a <=( a13791a  and  a13786a );
 a13795a <=( (not A168)  and  (not A169) );
 a13798a <=( A166  and  A167 );
 a13799a <=( a13798a  and  a13795a );
 a13802a <=( A233  and  A202 );
 a13806a <=( A267  and  A265 );
 a13807a <=( A234  and  a13806a );
 a13808a <=( a13807a  and  a13802a );
 a13811a <=( (not A168)  and  (not A169) );
 a13814a <=( A166  and  A167 );
 a13815a <=( a13814a  and  a13811a );
 a13818a <=( A233  and  A202 );
 a13822a <=( A267  and  A266 );
 a13823a <=( A234  and  a13822a );
 a13824a <=( a13823a  and  a13818a );
 a13827a <=( (not A168)  and  (not A169) );
 a13830a <=( A166  and  A167 );
 a13831a <=( a13830a  and  a13827a );
 a13834a <=( (not A232)  and  A202 );
 a13838a <=( A301  and  A236 );
 a13839a <=( A233  and  a13838a );
 a13840a <=( a13839a  and  a13834a );
 a13843a <=( (not A168)  and  (not A169) );
 a13846a <=( A166  and  A167 );
 a13847a <=( a13846a  and  a13843a );
 a13850a <=( (not A232)  and  A202 );
 a13854a <=( A268  and  A236 );
 a13855a <=( A233  and  a13854a );
 a13856a <=( a13855a  and  a13850a );
 a13859a <=( (not A168)  and  (not A169) );
 a13862a <=( A166  and  A167 );
 a13863a <=( a13862a  and  a13859a );
 a13866a <=( A232  and  A202 );
 a13870a <=( A301  and  A236 );
 a13871a <=( (not A233)  and  a13870a );
 a13872a <=( a13871a  and  a13866a );
 a13875a <=( (not A168)  and  (not A169) );
 a13878a <=( A166  and  A167 );
 a13879a <=( a13878a  and  a13875a );
 a13882a <=( A232  and  A202 );
 a13886a <=( A268  and  A236 );
 a13887a <=( (not A233)  and  a13886a );
 a13888a <=( a13887a  and  a13882a );
 a13891a <=( (not A168)  and  (not A169) );
 a13894a <=( A166  and  A167 );
 a13895a <=( a13894a  and  a13891a );
 a13898a <=( A201  and  A199 );
 a13902a <=( A300  and  A299 );
 a13903a <=( A235  and  a13902a );
 a13904a <=( a13903a  and  a13898a );
 a13907a <=( (not A168)  and  (not A169) );
 a13910a <=( A166  and  A167 );
 a13911a <=( a13910a  and  a13907a );
 a13914a <=( A201  and  A199 );
 a13918a <=( A300  and  A298 );
 a13919a <=( A235  and  a13918a );
 a13920a <=( a13919a  and  a13914a );
 a13923a <=( (not A168)  and  (not A169) );
 a13926a <=( A166  and  A167 );
 a13927a <=( a13926a  and  a13923a );
 a13930a <=( A201  and  A199 );
 a13934a <=( A267  and  A265 );
 a13935a <=( A235  and  a13934a );
 a13936a <=( a13935a  and  a13930a );
 a13939a <=( (not A168)  and  (not A169) );
 a13942a <=( A166  and  A167 );
 a13943a <=( a13942a  and  a13939a );
 a13946a <=( A201  and  A199 );
 a13950a <=( A267  and  A266 );
 a13951a <=( A235  and  a13950a );
 a13952a <=( a13951a  and  a13946a );
 a13955a <=( (not A168)  and  (not A169) );
 a13958a <=( A166  and  A167 );
 a13959a <=( a13958a  and  a13955a );
 a13962a <=( A201  and  A199 );
 a13966a <=( A301  and  A234 );
 a13967a <=( A232  and  a13966a );
 a13968a <=( a13967a  and  a13962a );
 a13971a <=( (not A168)  and  (not A169) );
 a13974a <=( A166  and  A167 );
 a13975a <=( a13974a  and  a13971a );
 a13978a <=( A201  and  A199 );
 a13982a <=( A268  and  A234 );
 a13983a <=( A232  and  a13982a );
 a13984a <=( a13983a  and  a13978a );
 a13987a <=( (not A168)  and  (not A169) );
 a13990a <=( A166  and  A167 );
 a13991a <=( a13990a  and  a13987a );
 a13994a <=( A201  and  A199 );
 a13998a <=( A301  and  A234 );
 a13999a <=( A233  and  a13998a );
 a14000a <=( a13999a  and  a13994a );
 a14003a <=( (not A168)  and  (not A169) );
 a14006a <=( A166  and  A167 );
 a14007a <=( a14006a  and  a14003a );
 a14010a <=( A201  and  A199 );
 a14014a <=( A268  and  A234 );
 a14015a <=( A233  and  a14014a );
 a14016a <=( a14015a  and  a14010a );
 a14019a <=( (not A168)  and  (not A169) );
 a14022a <=( A166  and  A167 );
 a14023a <=( a14022a  and  a14019a );
 a14026a <=( A201  and  A200 );
 a14030a <=( A300  and  A299 );
 a14031a <=( A235  and  a14030a );
 a14032a <=( a14031a  and  a14026a );
 a14035a <=( (not A168)  and  (not A169) );
 a14038a <=( A166  and  A167 );
 a14039a <=( a14038a  and  a14035a );
 a14042a <=( A201  and  A200 );
 a14046a <=( A300  and  A298 );
 a14047a <=( A235  and  a14046a );
 a14048a <=( a14047a  and  a14042a );
 a14051a <=( (not A168)  and  (not A169) );
 a14054a <=( A166  and  A167 );
 a14055a <=( a14054a  and  a14051a );
 a14058a <=( A201  and  A200 );
 a14062a <=( A267  and  A265 );
 a14063a <=( A235  and  a14062a );
 a14064a <=( a14063a  and  a14058a );
 a14067a <=( (not A168)  and  (not A169) );
 a14070a <=( A166  and  A167 );
 a14071a <=( a14070a  and  a14067a );
 a14074a <=( A201  and  A200 );
 a14078a <=( A267  and  A266 );
 a14079a <=( A235  and  a14078a );
 a14080a <=( a14079a  and  a14074a );
 a14083a <=( (not A168)  and  (not A169) );
 a14086a <=( A166  and  A167 );
 a14087a <=( a14086a  and  a14083a );
 a14090a <=( A201  and  A200 );
 a14094a <=( A301  and  A234 );
 a14095a <=( A232  and  a14094a );
 a14096a <=( a14095a  and  a14090a );
 a14099a <=( (not A168)  and  (not A169) );
 a14102a <=( A166  and  A167 );
 a14103a <=( a14102a  and  a14099a );
 a14106a <=( A201  and  A200 );
 a14110a <=( A268  and  A234 );
 a14111a <=( A232  and  a14110a );
 a14112a <=( a14111a  and  a14106a );
 a14115a <=( (not A168)  and  (not A169) );
 a14118a <=( A166  and  A167 );
 a14119a <=( a14118a  and  a14115a );
 a14122a <=( A201  and  A200 );
 a14126a <=( A301  and  A234 );
 a14127a <=( A233  and  a14126a );
 a14128a <=( a14127a  and  a14122a );
 a14131a <=( (not A168)  and  (not A169) );
 a14134a <=( A166  and  A167 );
 a14135a <=( a14134a  and  a14131a );
 a14138a <=( A201  and  A200 );
 a14142a <=( A268  and  A234 );
 a14143a <=( A233  and  a14142a );
 a14144a <=( a14143a  and  a14138a );
 a14147a <=( (not A168)  and  (not A169) );
 a14150a <=( A166  and  A167 );
 a14151a <=( a14150a  and  a14147a );
 a14154a <=( A200  and  (not A199) );
 a14158a <=( A301  and  A235 );
 a14159a <=( A203  and  a14158a );
 a14160a <=( a14159a  and  a14154a );
 a14163a <=( (not A168)  and  (not A169) );
 a14166a <=( A166  and  A167 );
 a14167a <=( a14166a  and  a14163a );
 a14170a <=( A200  and  (not A199) );
 a14174a <=( A268  and  A235 );
 a14175a <=( A203  and  a14174a );
 a14176a <=( a14175a  and  a14170a );
 a14179a <=( (not A168)  and  (not A169) );
 a14182a <=( A166  and  A167 );
 a14183a <=( a14182a  and  a14179a );
 a14186a <=( (not A200)  and  A199 );
 a14190a <=( A301  and  A235 );
 a14191a <=( A203  and  a14190a );
 a14192a <=( a14191a  and  a14186a );
 a14195a <=( (not A168)  and  (not A169) );
 a14198a <=( A166  and  A167 );
 a14199a <=( a14198a  and  a14195a );
 a14202a <=( (not A200)  and  A199 );
 a14206a <=( A268  and  A235 );
 a14207a <=( A203  and  a14206a );
 a14208a <=( a14207a  and  a14202a );
 a14211a <=( (not A169)  and  (not A170) );
 a14214a <=( A202  and  (not A168) );
 a14215a <=( a14214a  and  a14211a );
 a14218a <=( A234  and  A232 );
 a14222a <=( A302  and  (not A299) );
 a14223a <=( A298  and  a14222a );
 a14224a <=( a14223a  and  a14218a );
 a14227a <=( (not A169)  and  (not A170) );
 a14230a <=( A202  and  (not A168) );
 a14231a <=( a14230a  and  a14227a );
 a14234a <=( A234  and  A232 );
 a14238a <=( A302  and  A299 );
 a14239a <=( (not A298)  and  a14238a );
 a14240a <=( a14239a  and  a14234a );
 a14243a <=( (not A169)  and  (not A170) );
 a14246a <=( A202  and  (not A168) );
 a14247a <=( a14246a  and  a14243a );
 a14250a <=( A234  and  A232 );
 a14254a <=( A269  and  A266 );
 a14255a <=( (not A265)  and  a14254a );
 a14256a <=( a14255a  and  a14250a );
 a14259a <=( (not A169)  and  (not A170) );
 a14262a <=( A202  and  (not A168) );
 a14263a <=( a14262a  and  a14259a );
 a14266a <=( A234  and  A232 );
 a14270a <=( A269  and  (not A266) );
 a14271a <=( A265  and  a14270a );
 a14272a <=( a14271a  and  a14266a );
 a14275a <=( (not A169)  and  (not A170) );
 a14278a <=( A202  and  (not A168) );
 a14279a <=( a14278a  and  a14275a );
 a14282a <=( A234  and  A233 );
 a14286a <=( A302  and  (not A299) );
 a14287a <=( A298  and  a14286a );
 a14288a <=( a14287a  and  a14282a );
 a14291a <=( (not A169)  and  (not A170) );
 a14294a <=( A202  and  (not A168) );
 a14295a <=( a14294a  and  a14291a );
 a14298a <=( A234  and  A233 );
 a14302a <=( A302  and  A299 );
 a14303a <=( (not A298)  and  a14302a );
 a14304a <=( a14303a  and  a14298a );
 a14307a <=( (not A169)  and  (not A170) );
 a14310a <=( A202  and  (not A168) );
 a14311a <=( a14310a  and  a14307a );
 a14314a <=( A234  and  A233 );
 a14318a <=( A269  and  A266 );
 a14319a <=( (not A265)  and  a14318a );
 a14320a <=( a14319a  and  a14314a );
 a14323a <=( (not A169)  and  (not A170) );
 a14326a <=( A202  and  (not A168) );
 a14327a <=( a14326a  and  a14323a );
 a14330a <=( A234  and  A233 );
 a14334a <=( A269  and  (not A266) );
 a14335a <=( A265  and  a14334a );
 a14336a <=( a14335a  and  a14330a );
 a14339a <=( (not A169)  and  (not A170) );
 a14342a <=( A202  and  (not A168) );
 a14343a <=( a14342a  and  a14339a );
 a14346a <=( A233  and  (not A232) );
 a14350a <=( A300  and  A299 );
 a14351a <=( A236  and  a14350a );
 a14352a <=( a14351a  and  a14346a );
 a14355a <=( (not A169)  and  (not A170) );
 a14358a <=( A202  and  (not A168) );
 a14359a <=( a14358a  and  a14355a );
 a14362a <=( A233  and  (not A232) );
 a14366a <=( A300  and  A298 );
 a14367a <=( A236  and  a14366a );
 a14368a <=( a14367a  and  a14362a );
 a14371a <=( (not A169)  and  (not A170) );
 a14374a <=( A202  and  (not A168) );
 a14375a <=( a14374a  and  a14371a );
 a14378a <=( A233  and  (not A232) );
 a14382a <=( A267  and  A265 );
 a14383a <=( A236  and  a14382a );
 a14384a <=( a14383a  and  a14378a );
 a14387a <=( (not A169)  and  (not A170) );
 a14390a <=( A202  and  (not A168) );
 a14391a <=( a14390a  and  a14387a );
 a14394a <=( A233  and  (not A232) );
 a14398a <=( A267  and  A266 );
 a14399a <=( A236  and  a14398a );
 a14400a <=( a14399a  and  a14394a );
 a14403a <=( (not A169)  and  (not A170) );
 a14406a <=( A202  and  (not A168) );
 a14407a <=( a14406a  and  a14403a );
 a14410a <=( (not A233)  and  A232 );
 a14414a <=( A300  and  A299 );
 a14415a <=( A236  and  a14414a );
 a14416a <=( a14415a  and  a14410a );
 a14419a <=( (not A169)  and  (not A170) );
 a14422a <=( A202  and  (not A168) );
 a14423a <=( a14422a  and  a14419a );
 a14426a <=( (not A233)  and  A232 );
 a14430a <=( A300  and  A298 );
 a14431a <=( A236  and  a14430a );
 a14432a <=( a14431a  and  a14426a );
 a14435a <=( (not A169)  and  (not A170) );
 a14438a <=( A202  and  (not A168) );
 a14439a <=( a14438a  and  a14435a );
 a14442a <=( (not A233)  and  A232 );
 a14446a <=( A267  and  A265 );
 a14447a <=( A236  and  a14446a );
 a14448a <=( a14447a  and  a14442a );
 a14451a <=( (not A169)  and  (not A170) );
 a14454a <=( A202  and  (not A168) );
 a14455a <=( a14454a  and  a14451a );
 a14458a <=( (not A233)  and  A232 );
 a14462a <=( A267  and  A266 );
 a14463a <=( A236  and  a14462a );
 a14464a <=( a14463a  and  a14458a );
 a14467a <=( (not A169)  and  (not A170) );
 a14470a <=( A199  and  (not A168) );
 a14471a <=( a14470a  and  a14467a );
 a14474a <=( A235  and  A201 );
 a14478a <=( A302  and  (not A299) );
 a14479a <=( A298  and  a14478a );
 a14480a <=( a14479a  and  a14474a );
 a14483a <=( (not A169)  and  (not A170) );
 a14486a <=( A199  and  (not A168) );
 a14487a <=( a14486a  and  a14483a );
 a14490a <=( A235  and  A201 );
 a14494a <=( A302  and  A299 );
 a14495a <=( (not A298)  and  a14494a );
 a14496a <=( a14495a  and  a14490a );
 a14499a <=( (not A169)  and  (not A170) );
 a14502a <=( A199  and  (not A168) );
 a14503a <=( a14502a  and  a14499a );
 a14506a <=( A235  and  A201 );
 a14510a <=( A269  and  A266 );
 a14511a <=( (not A265)  and  a14510a );
 a14512a <=( a14511a  and  a14506a );
 a14515a <=( (not A169)  and  (not A170) );
 a14518a <=( A199  and  (not A168) );
 a14519a <=( a14518a  and  a14515a );
 a14522a <=( A235  and  A201 );
 a14526a <=( A269  and  (not A266) );
 a14527a <=( A265  and  a14526a );
 a14528a <=( a14527a  and  a14522a );
 a14531a <=( (not A169)  and  (not A170) );
 a14534a <=( A199  and  (not A168) );
 a14535a <=( a14534a  and  a14531a );
 a14538a <=( A232  and  A201 );
 a14542a <=( A300  and  A299 );
 a14543a <=( A234  and  a14542a );
 a14544a <=( a14543a  and  a14538a );
 a14547a <=( (not A169)  and  (not A170) );
 a14550a <=( A199  and  (not A168) );
 a14551a <=( a14550a  and  a14547a );
 a14554a <=( A232  and  A201 );
 a14558a <=( A300  and  A298 );
 a14559a <=( A234  and  a14558a );
 a14560a <=( a14559a  and  a14554a );
 a14563a <=( (not A169)  and  (not A170) );
 a14566a <=( A199  and  (not A168) );
 a14567a <=( a14566a  and  a14563a );
 a14570a <=( A232  and  A201 );
 a14574a <=( A267  and  A265 );
 a14575a <=( A234  and  a14574a );
 a14576a <=( a14575a  and  a14570a );
 a14579a <=( (not A169)  and  (not A170) );
 a14582a <=( A199  and  (not A168) );
 a14583a <=( a14582a  and  a14579a );
 a14586a <=( A232  and  A201 );
 a14590a <=( A267  and  A266 );
 a14591a <=( A234  and  a14590a );
 a14592a <=( a14591a  and  a14586a );
 a14595a <=( (not A169)  and  (not A170) );
 a14598a <=( A199  and  (not A168) );
 a14599a <=( a14598a  and  a14595a );
 a14602a <=( A233  and  A201 );
 a14606a <=( A300  and  A299 );
 a14607a <=( A234  and  a14606a );
 a14608a <=( a14607a  and  a14602a );
 a14611a <=( (not A169)  and  (not A170) );
 a14614a <=( A199  and  (not A168) );
 a14615a <=( a14614a  and  a14611a );
 a14618a <=( A233  and  A201 );
 a14622a <=( A300  and  A298 );
 a14623a <=( A234  and  a14622a );
 a14624a <=( a14623a  and  a14618a );
 a14627a <=( (not A169)  and  (not A170) );
 a14630a <=( A199  and  (not A168) );
 a14631a <=( a14630a  and  a14627a );
 a14634a <=( A233  and  A201 );
 a14638a <=( A267  and  A265 );
 a14639a <=( A234  and  a14638a );
 a14640a <=( a14639a  and  a14634a );
 a14643a <=( (not A169)  and  (not A170) );
 a14646a <=( A199  and  (not A168) );
 a14647a <=( a14646a  and  a14643a );
 a14650a <=( A233  and  A201 );
 a14654a <=( A267  and  A266 );
 a14655a <=( A234  and  a14654a );
 a14656a <=( a14655a  and  a14650a );
 a14659a <=( (not A169)  and  (not A170) );
 a14662a <=( A199  and  (not A168) );
 a14663a <=( a14662a  and  a14659a );
 a14666a <=( (not A232)  and  A201 );
 a14670a <=( A301  and  A236 );
 a14671a <=( A233  and  a14670a );
 a14672a <=( a14671a  and  a14666a );
 a14675a <=( (not A169)  and  (not A170) );
 a14678a <=( A199  and  (not A168) );
 a14679a <=( a14678a  and  a14675a );
 a14682a <=( (not A232)  and  A201 );
 a14686a <=( A268  and  A236 );
 a14687a <=( A233  and  a14686a );
 a14688a <=( a14687a  and  a14682a );
 a14691a <=( (not A169)  and  (not A170) );
 a14694a <=( A199  and  (not A168) );
 a14695a <=( a14694a  and  a14691a );
 a14698a <=( A232  and  A201 );
 a14702a <=( A301  and  A236 );
 a14703a <=( (not A233)  and  a14702a );
 a14704a <=( a14703a  and  a14698a );
 a14707a <=( (not A169)  and  (not A170) );
 a14710a <=( A199  and  (not A168) );
 a14711a <=( a14710a  and  a14707a );
 a14714a <=( A232  and  A201 );
 a14718a <=( A268  and  A236 );
 a14719a <=( (not A233)  and  a14718a );
 a14720a <=( a14719a  and  a14714a );
 a14723a <=( (not A169)  and  (not A170) );
 a14726a <=( A200  and  (not A168) );
 a14727a <=( a14726a  and  a14723a );
 a14730a <=( A235  and  A201 );
 a14734a <=( A302  and  (not A299) );
 a14735a <=( A298  and  a14734a );
 a14736a <=( a14735a  and  a14730a );
 a14739a <=( (not A169)  and  (not A170) );
 a14742a <=( A200  and  (not A168) );
 a14743a <=( a14742a  and  a14739a );
 a14746a <=( A235  and  A201 );
 a14750a <=( A302  and  A299 );
 a14751a <=( (not A298)  and  a14750a );
 a14752a <=( a14751a  and  a14746a );
 a14755a <=( (not A169)  and  (not A170) );
 a14758a <=( A200  and  (not A168) );
 a14759a <=( a14758a  and  a14755a );
 a14762a <=( A235  and  A201 );
 a14766a <=( A269  and  A266 );
 a14767a <=( (not A265)  and  a14766a );
 a14768a <=( a14767a  and  a14762a );
 a14771a <=( (not A169)  and  (not A170) );
 a14774a <=( A200  and  (not A168) );
 a14775a <=( a14774a  and  a14771a );
 a14778a <=( A235  and  A201 );
 a14782a <=( A269  and  (not A266) );
 a14783a <=( A265  and  a14782a );
 a14784a <=( a14783a  and  a14778a );
 a14787a <=( (not A169)  and  (not A170) );
 a14790a <=( A200  and  (not A168) );
 a14791a <=( a14790a  and  a14787a );
 a14794a <=( A232  and  A201 );
 a14798a <=( A300  and  A299 );
 a14799a <=( A234  and  a14798a );
 a14800a <=( a14799a  and  a14794a );
 a14803a <=( (not A169)  and  (not A170) );
 a14806a <=( A200  and  (not A168) );
 a14807a <=( a14806a  and  a14803a );
 a14810a <=( A232  and  A201 );
 a14814a <=( A300  and  A298 );
 a14815a <=( A234  and  a14814a );
 a14816a <=( a14815a  and  a14810a );
 a14819a <=( (not A169)  and  (not A170) );
 a14822a <=( A200  and  (not A168) );
 a14823a <=( a14822a  and  a14819a );
 a14826a <=( A232  and  A201 );
 a14830a <=( A267  and  A265 );
 a14831a <=( A234  and  a14830a );
 a14832a <=( a14831a  and  a14826a );
 a14835a <=( (not A169)  and  (not A170) );
 a14838a <=( A200  and  (not A168) );
 a14839a <=( a14838a  and  a14835a );
 a14842a <=( A232  and  A201 );
 a14846a <=( A267  and  A266 );
 a14847a <=( A234  and  a14846a );
 a14848a <=( a14847a  and  a14842a );
 a14851a <=( (not A169)  and  (not A170) );
 a14854a <=( A200  and  (not A168) );
 a14855a <=( a14854a  and  a14851a );
 a14858a <=( A233  and  A201 );
 a14862a <=( A300  and  A299 );
 a14863a <=( A234  and  a14862a );
 a14864a <=( a14863a  and  a14858a );
 a14867a <=( (not A169)  and  (not A170) );
 a14870a <=( A200  and  (not A168) );
 a14871a <=( a14870a  and  a14867a );
 a14874a <=( A233  and  A201 );
 a14878a <=( A300  and  A298 );
 a14879a <=( A234  and  a14878a );
 a14880a <=( a14879a  and  a14874a );
 a14883a <=( (not A169)  and  (not A170) );
 a14886a <=( A200  and  (not A168) );
 a14887a <=( a14886a  and  a14883a );
 a14890a <=( A233  and  A201 );
 a14894a <=( A267  and  A265 );
 a14895a <=( A234  and  a14894a );
 a14896a <=( a14895a  and  a14890a );
 a14899a <=( (not A169)  and  (not A170) );
 a14902a <=( A200  and  (not A168) );
 a14903a <=( a14902a  and  a14899a );
 a14906a <=( A233  and  A201 );
 a14910a <=( A267  and  A266 );
 a14911a <=( A234  and  a14910a );
 a14912a <=( a14911a  and  a14906a );
 a14915a <=( (not A169)  and  (not A170) );
 a14918a <=( A200  and  (not A168) );
 a14919a <=( a14918a  and  a14915a );
 a14922a <=( (not A232)  and  A201 );
 a14926a <=( A301  and  A236 );
 a14927a <=( A233  and  a14926a );
 a14928a <=( a14927a  and  a14922a );
 a14931a <=( (not A169)  and  (not A170) );
 a14934a <=( A200  and  (not A168) );
 a14935a <=( a14934a  and  a14931a );
 a14938a <=( (not A232)  and  A201 );
 a14942a <=( A268  and  A236 );
 a14943a <=( A233  and  a14942a );
 a14944a <=( a14943a  and  a14938a );
 a14947a <=( (not A169)  and  (not A170) );
 a14950a <=( A200  and  (not A168) );
 a14951a <=( a14950a  and  a14947a );
 a14954a <=( A232  and  A201 );
 a14958a <=( A301  and  A236 );
 a14959a <=( (not A233)  and  a14958a );
 a14960a <=( a14959a  and  a14954a );
 a14963a <=( (not A169)  and  (not A170) );
 a14966a <=( A200  and  (not A168) );
 a14967a <=( a14966a  and  a14963a );
 a14970a <=( A232  and  A201 );
 a14974a <=( A268  and  A236 );
 a14975a <=( (not A233)  and  a14974a );
 a14976a <=( a14975a  and  a14970a );
 a14979a <=( (not A169)  and  (not A170) );
 a14982a <=( (not A199)  and  (not A168) );
 a14983a <=( a14982a  and  a14979a );
 a14986a <=( A203  and  A200 );
 a14990a <=( A300  and  A299 );
 a14991a <=( A235  and  a14990a );
 a14992a <=( a14991a  and  a14986a );
 a14995a <=( (not A169)  and  (not A170) );
 a14998a <=( (not A199)  and  (not A168) );
 a14999a <=( a14998a  and  a14995a );
 a15002a <=( A203  and  A200 );
 a15006a <=( A300  and  A298 );
 a15007a <=( A235  and  a15006a );
 a15008a <=( a15007a  and  a15002a );
 a15011a <=( (not A169)  and  (not A170) );
 a15014a <=( (not A199)  and  (not A168) );
 a15015a <=( a15014a  and  a15011a );
 a15018a <=( A203  and  A200 );
 a15022a <=( A267  and  A265 );
 a15023a <=( A235  and  a15022a );
 a15024a <=( a15023a  and  a15018a );
 a15027a <=( (not A169)  and  (not A170) );
 a15030a <=( (not A199)  and  (not A168) );
 a15031a <=( a15030a  and  a15027a );
 a15034a <=( A203  and  A200 );
 a15038a <=( A267  and  A266 );
 a15039a <=( A235  and  a15038a );
 a15040a <=( a15039a  and  a15034a );
 a15043a <=( (not A169)  and  (not A170) );
 a15046a <=( (not A199)  and  (not A168) );
 a15047a <=( a15046a  and  a15043a );
 a15050a <=( A203  and  A200 );
 a15054a <=( A301  and  A234 );
 a15055a <=( A232  and  a15054a );
 a15056a <=( a15055a  and  a15050a );
 a15059a <=( (not A169)  and  (not A170) );
 a15062a <=( (not A199)  and  (not A168) );
 a15063a <=( a15062a  and  a15059a );
 a15066a <=( A203  and  A200 );
 a15070a <=( A268  and  A234 );
 a15071a <=( A232  and  a15070a );
 a15072a <=( a15071a  and  a15066a );
 a15075a <=( (not A169)  and  (not A170) );
 a15078a <=( (not A199)  and  (not A168) );
 a15079a <=( a15078a  and  a15075a );
 a15082a <=( A203  and  A200 );
 a15086a <=( A301  and  A234 );
 a15087a <=( A233  and  a15086a );
 a15088a <=( a15087a  and  a15082a );
 a15091a <=( (not A169)  and  (not A170) );
 a15094a <=( (not A199)  and  (not A168) );
 a15095a <=( a15094a  and  a15091a );
 a15098a <=( A203  and  A200 );
 a15102a <=( A268  and  A234 );
 a15103a <=( A233  and  a15102a );
 a15104a <=( a15103a  and  a15098a );
 a15107a <=( (not A169)  and  (not A170) );
 a15110a <=( A199  and  (not A168) );
 a15111a <=( a15110a  and  a15107a );
 a15114a <=( A203  and  (not A200) );
 a15118a <=( A300  and  A299 );
 a15119a <=( A235  and  a15118a );
 a15120a <=( a15119a  and  a15114a );
 a15123a <=( (not A169)  and  (not A170) );
 a15126a <=( A199  and  (not A168) );
 a15127a <=( a15126a  and  a15123a );
 a15130a <=( A203  and  (not A200) );
 a15134a <=( A300  and  A298 );
 a15135a <=( A235  and  a15134a );
 a15136a <=( a15135a  and  a15130a );
 a15139a <=( (not A169)  and  (not A170) );
 a15142a <=( A199  and  (not A168) );
 a15143a <=( a15142a  and  a15139a );
 a15146a <=( A203  and  (not A200) );
 a15150a <=( A267  and  A265 );
 a15151a <=( A235  and  a15150a );
 a15152a <=( a15151a  and  a15146a );
 a15155a <=( (not A169)  and  (not A170) );
 a15158a <=( A199  and  (not A168) );
 a15159a <=( a15158a  and  a15155a );
 a15162a <=( A203  and  (not A200) );
 a15166a <=( A267  and  A266 );
 a15167a <=( A235  and  a15166a );
 a15168a <=( a15167a  and  a15162a );
 a15171a <=( (not A169)  and  (not A170) );
 a15174a <=( A199  and  (not A168) );
 a15175a <=( a15174a  and  a15171a );
 a15178a <=( A203  and  (not A200) );
 a15182a <=( A301  and  A234 );
 a15183a <=( A232  and  a15182a );
 a15184a <=( a15183a  and  a15178a );
 a15187a <=( (not A169)  and  (not A170) );
 a15190a <=( A199  and  (not A168) );
 a15191a <=( a15190a  and  a15187a );
 a15194a <=( A203  and  (not A200) );
 a15198a <=( A268  and  A234 );
 a15199a <=( A232  and  a15198a );
 a15200a <=( a15199a  and  a15194a );
 a15203a <=( (not A169)  and  (not A170) );
 a15206a <=( A199  and  (not A168) );
 a15207a <=( a15206a  and  a15203a );
 a15210a <=( A203  and  (not A200) );
 a15214a <=( A301  and  A234 );
 a15215a <=( A233  and  a15214a );
 a15216a <=( a15215a  and  a15210a );
 a15219a <=( (not A169)  and  (not A170) );
 a15222a <=( A199  and  (not A168) );
 a15223a <=( a15222a  and  a15219a );
 a15226a <=( A203  and  (not A200) );
 a15230a <=( A268  and  A234 );
 a15231a <=( A233  and  a15230a );
 a15232a <=( a15231a  and  a15226a );
 a15235a <=( A166  and  A168 );
 a15239a <=( (not A203)  and  (not A202) );
 a15240a <=( (not A201)  and  a15239a );
 a15241a <=( a15240a  and  a15235a );
 a15244a <=( A234  and  A232 );
 a15248a <=( A302  and  (not A299) );
 a15249a <=( A298  and  a15248a );
 a15250a <=( a15249a  and  a15244a );
 a15253a <=( A166  and  A168 );
 a15257a <=( (not A203)  and  (not A202) );
 a15258a <=( (not A201)  and  a15257a );
 a15259a <=( a15258a  and  a15253a );
 a15262a <=( A234  and  A232 );
 a15266a <=( A302  and  A299 );
 a15267a <=( (not A298)  and  a15266a );
 a15268a <=( a15267a  and  a15262a );
 a15271a <=( A166  and  A168 );
 a15275a <=( (not A203)  and  (not A202) );
 a15276a <=( (not A201)  and  a15275a );
 a15277a <=( a15276a  and  a15271a );
 a15280a <=( A234  and  A232 );
 a15284a <=( A269  and  A266 );
 a15285a <=( (not A265)  and  a15284a );
 a15286a <=( a15285a  and  a15280a );
 a15289a <=( A166  and  A168 );
 a15293a <=( (not A203)  and  (not A202) );
 a15294a <=( (not A201)  and  a15293a );
 a15295a <=( a15294a  and  a15289a );
 a15298a <=( A234  and  A232 );
 a15302a <=( A269  and  (not A266) );
 a15303a <=( A265  and  a15302a );
 a15304a <=( a15303a  and  a15298a );
 a15307a <=( A166  and  A168 );
 a15311a <=( (not A203)  and  (not A202) );
 a15312a <=( (not A201)  and  a15311a );
 a15313a <=( a15312a  and  a15307a );
 a15316a <=( A234  and  A233 );
 a15320a <=( A302  and  (not A299) );
 a15321a <=( A298  and  a15320a );
 a15322a <=( a15321a  and  a15316a );
 a15325a <=( A166  and  A168 );
 a15329a <=( (not A203)  and  (not A202) );
 a15330a <=( (not A201)  and  a15329a );
 a15331a <=( a15330a  and  a15325a );
 a15334a <=( A234  and  A233 );
 a15338a <=( A302  and  A299 );
 a15339a <=( (not A298)  and  a15338a );
 a15340a <=( a15339a  and  a15334a );
 a15343a <=( A166  and  A168 );
 a15347a <=( (not A203)  and  (not A202) );
 a15348a <=( (not A201)  and  a15347a );
 a15349a <=( a15348a  and  a15343a );
 a15352a <=( A234  and  A233 );
 a15356a <=( A269  and  A266 );
 a15357a <=( (not A265)  and  a15356a );
 a15358a <=( a15357a  and  a15352a );
 a15361a <=( A166  and  A168 );
 a15365a <=( (not A203)  and  (not A202) );
 a15366a <=( (not A201)  and  a15365a );
 a15367a <=( a15366a  and  a15361a );
 a15370a <=( A234  and  A233 );
 a15374a <=( A269  and  (not A266) );
 a15375a <=( A265  and  a15374a );
 a15376a <=( a15375a  and  a15370a );
 a15379a <=( A166  and  A168 );
 a15383a <=( (not A203)  and  (not A202) );
 a15384a <=( (not A201)  and  a15383a );
 a15385a <=( a15384a  and  a15379a );
 a15388a <=( A233  and  (not A232) );
 a15392a <=( A300  and  A299 );
 a15393a <=( A236  and  a15392a );
 a15394a <=( a15393a  and  a15388a );
 a15397a <=( A166  and  A168 );
 a15401a <=( (not A203)  and  (not A202) );
 a15402a <=( (not A201)  and  a15401a );
 a15403a <=( a15402a  and  a15397a );
 a15406a <=( A233  and  (not A232) );
 a15410a <=( A300  and  A298 );
 a15411a <=( A236  and  a15410a );
 a15412a <=( a15411a  and  a15406a );
 a15415a <=( A166  and  A168 );
 a15419a <=( (not A203)  and  (not A202) );
 a15420a <=( (not A201)  and  a15419a );
 a15421a <=( a15420a  and  a15415a );
 a15424a <=( A233  and  (not A232) );
 a15428a <=( A267  and  A265 );
 a15429a <=( A236  and  a15428a );
 a15430a <=( a15429a  and  a15424a );
 a15433a <=( A166  and  A168 );
 a15437a <=( (not A203)  and  (not A202) );
 a15438a <=( (not A201)  and  a15437a );
 a15439a <=( a15438a  and  a15433a );
 a15442a <=( A233  and  (not A232) );
 a15446a <=( A267  and  A266 );
 a15447a <=( A236  and  a15446a );
 a15448a <=( a15447a  and  a15442a );
 a15451a <=( A166  and  A168 );
 a15455a <=( (not A203)  and  (not A202) );
 a15456a <=( (not A201)  and  a15455a );
 a15457a <=( a15456a  and  a15451a );
 a15460a <=( (not A233)  and  A232 );
 a15464a <=( A300  and  A299 );
 a15465a <=( A236  and  a15464a );
 a15466a <=( a15465a  and  a15460a );
 a15469a <=( A166  and  A168 );
 a15473a <=( (not A203)  and  (not A202) );
 a15474a <=( (not A201)  and  a15473a );
 a15475a <=( a15474a  and  a15469a );
 a15478a <=( (not A233)  and  A232 );
 a15482a <=( A300  and  A298 );
 a15483a <=( A236  and  a15482a );
 a15484a <=( a15483a  and  a15478a );
 a15487a <=( A166  and  A168 );
 a15491a <=( (not A203)  and  (not A202) );
 a15492a <=( (not A201)  and  a15491a );
 a15493a <=( a15492a  and  a15487a );
 a15496a <=( (not A233)  and  A232 );
 a15500a <=( A267  and  A265 );
 a15501a <=( A236  and  a15500a );
 a15502a <=( a15501a  and  a15496a );
 a15505a <=( A166  and  A168 );
 a15509a <=( (not A203)  and  (not A202) );
 a15510a <=( (not A201)  and  a15509a );
 a15511a <=( a15510a  and  a15505a );
 a15514a <=( (not A233)  and  A232 );
 a15518a <=( A267  and  A266 );
 a15519a <=( A236  and  a15518a );
 a15520a <=( a15519a  and  a15514a );
 a15523a <=( A166  and  A168 );
 a15527a <=( (not A201)  and  A200 );
 a15528a <=( A199  and  a15527a );
 a15529a <=( a15528a  and  a15523a );
 a15532a <=( A235  and  (not A202) );
 a15536a <=( A302  and  (not A299) );
 a15537a <=( A298  and  a15536a );
 a15538a <=( a15537a  and  a15532a );
 a15541a <=( A166  and  A168 );
 a15545a <=( (not A201)  and  A200 );
 a15546a <=( A199  and  a15545a );
 a15547a <=( a15546a  and  a15541a );
 a15550a <=( A235  and  (not A202) );
 a15554a <=( A302  and  A299 );
 a15555a <=( (not A298)  and  a15554a );
 a15556a <=( a15555a  and  a15550a );
 a15559a <=( A166  and  A168 );
 a15563a <=( (not A201)  and  A200 );
 a15564a <=( A199  and  a15563a );
 a15565a <=( a15564a  and  a15559a );
 a15568a <=( A235  and  (not A202) );
 a15572a <=( A269  and  A266 );
 a15573a <=( (not A265)  and  a15572a );
 a15574a <=( a15573a  and  a15568a );
 a15577a <=( A166  and  A168 );
 a15581a <=( (not A201)  and  A200 );
 a15582a <=( A199  and  a15581a );
 a15583a <=( a15582a  and  a15577a );
 a15586a <=( A235  and  (not A202) );
 a15590a <=( A269  and  (not A266) );
 a15591a <=( A265  and  a15590a );
 a15592a <=( a15591a  and  a15586a );
 a15595a <=( A166  and  A168 );
 a15599a <=( (not A201)  and  A200 );
 a15600a <=( A199  and  a15599a );
 a15601a <=( a15600a  and  a15595a );
 a15604a <=( A232  and  (not A202) );
 a15608a <=( A300  and  A299 );
 a15609a <=( A234  and  a15608a );
 a15610a <=( a15609a  and  a15604a );
 a15613a <=( A166  and  A168 );
 a15617a <=( (not A201)  and  A200 );
 a15618a <=( A199  and  a15617a );
 a15619a <=( a15618a  and  a15613a );
 a15622a <=( A232  and  (not A202) );
 a15626a <=( A300  and  A298 );
 a15627a <=( A234  and  a15626a );
 a15628a <=( a15627a  and  a15622a );
 a15631a <=( A166  and  A168 );
 a15635a <=( (not A201)  and  A200 );
 a15636a <=( A199  and  a15635a );
 a15637a <=( a15636a  and  a15631a );
 a15640a <=( A232  and  (not A202) );
 a15644a <=( A267  and  A265 );
 a15645a <=( A234  and  a15644a );
 a15646a <=( a15645a  and  a15640a );
 a15649a <=( A166  and  A168 );
 a15653a <=( (not A201)  and  A200 );
 a15654a <=( A199  and  a15653a );
 a15655a <=( a15654a  and  a15649a );
 a15658a <=( A232  and  (not A202) );
 a15662a <=( A267  and  A266 );
 a15663a <=( A234  and  a15662a );
 a15664a <=( a15663a  and  a15658a );
 a15667a <=( A166  and  A168 );
 a15671a <=( (not A201)  and  A200 );
 a15672a <=( A199  and  a15671a );
 a15673a <=( a15672a  and  a15667a );
 a15676a <=( A233  and  (not A202) );
 a15680a <=( A300  and  A299 );
 a15681a <=( A234  and  a15680a );
 a15682a <=( a15681a  and  a15676a );
 a15685a <=( A166  and  A168 );
 a15689a <=( (not A201)  and  A200 );
 a15690a <=( A199  and  a15689a );
 a15691a <=( a15690a  and  a15685a );
 a15694a <=( A233  and  (not A202) );
 a15698a <=( A300  and  A298 );
 a15699a <=( A234  and  a15698a );
 a15700a <=( a15699a  and  a15694a );
 a15703a <=( A166  and  A168 );
 a15707a <=( (not A201)  and  A200 );
 a15708a <=( A199  and  a15707a );
 a15709a <=( a15708a  and  a15703a );
 a15712a <=( A233  and  (not A202) );
 a15716a <=( A267  and  A265 );
 a15717a <=( A234  and  a15716a );
 a15718a <=( a15717a  and  a15712a );
 a15721a <=( A166  and  A168 );
 a15725a <=( (not A201)  and  A200 );
 a15726a <=( A199  and  a15725a );
 a15727a <=( a15726a  and  a15721a );
 a15730a <=( A233  and  (not A202) );
 a15734a <=( A267  and  A266 );
 a15735a <=( A234  and  a15734a );
 a15736a <=( a15735a  and  a15730a );
 a15739a <=( A166  and  A168 );
 a15743a <=( (not A201)  and  A200 );
 a15744a <=( A199  and  a15743a );
 a15745a <=( a15744a  and  a15739a );
 a15748a <=( (not A232)  and  (not A202) );
 a15752a <=( A301  and  A236 );
 a15753a <=( A233  and  a15752a );
 a15754a <=( a15753a  and  a15748a );
 a15757a <=( A166  and  A168 );
 a15761a <=( (not A201)  and  A200 );
 a15762a <=( A199  and  a15761a );
 a15763a <=( a15762a  and  a15757a );
 a15766a <=( (not A232)  and  (not A202) );
 a15770a <=( A268  and  A236 );
 a15771a <=( A233  and  a15770a );
 a15772a <=( a15771a  and  a15766a );
 a15775a <=( A166  and  A168 );
 a15779a <=( (not A201)  and  A200 );
 a15780a <=( A199  and  a15779a );
 a15781a <=( a15780a  and  a15775a );
 a15784a <=( A232  and  (not A202) );
 a15788a <=( A301  and  A236 );
 a15789a <=( (not A233)  and  a15788a );
 a15790a <=( a15789a  and  a15784a );
 a15793a <=( A166  and  A168 );
 a15797a <=( (not A201)  and  A200 );
 a15798a <=( A199  and  a15797a );
 a15799a <=( a15798a  and  a15793a );
 a15802a <=( A232  and  (not A202) );
 a15806a <=( A268  and  A236 );
 a15807a <=( (not A233)  and  a15806a );
 a15808a <=( a15807a  and  a15802a );
 a15811a <=( A166  and  A168 );
 a15815a <=( (not A202)  and  (not A200) );
 a15816a <=( (not A199)  and  a15815a );
 a15817a <=( a15816a  and  a15811a );
 a15820a <=( A234  and  A232 );
 a15824a <=( A302  and  (not A299) );
 a15825a <=( A298  and  a15824a );
 a15826a <=( a15825a  and  a15820a );
 a15829a <=( A166  and  A168 );
 a15833a <=( (not A202)  and  (not A200) );
 a15834a <=( (not A199)  and  a15833a );
 a15835a <=( a15834a  and  a15829a );
 a15838a <=( A234  and  A232 );
 a15842a <=( A302  and  A299 );
 a15843a <=( (not A298)  and  a15842a );
 a15844a <=( a15843a  and  a15838a );
 a15847a <=( A166  and  A168 );
 a15851a <=( (not A202)  and  (not A200) );
 a15852a <=( (not A199)  and  a15851a );
 a15853a <=( a15852a  and  a15847a );
 a15856a <=( A234  and  A232 );
 a15860a <=( A269  and  A266 );
 a15861a <=( (not A265)  and  a15860a );
 a15862a <=( a15861a  and  a15856a );
 a15865a <=( A166  and  A168 );
 a15869a <=( (not A202)  and  (not A200) );
 a15870a <=( (not A199)  and  a15869a );
 a15871a <=( a15870a  and  a15865a );
 a15874a <=( A234  and  A232 );
 a15878a <=( A269  and  (not A266) );
 a15879a <=( A265  and  a15878a );
 a15880a <=( a15879a  and  a15874a );
 a15883a <=( A166  and  A168 );
 a15887a <=( (not A202)  and  (not A200) );
 a15888a <=( (not A199)  and  a15887a );
 a15889a <=( a15888a  and  a15883a );
 a15892a <=( A234  and  A233 );
 a15896a <=( A302  and  (not A299) );
 a15897a <=( A298  and  a15896a );
 a15898a <=( a15897a  and  a15892a );
 a15901a <=( A166  and  A168 );
 a15905a <=( (not A202)  and  (not A200) );
 a15906a <=( (not A199)  and  a15905a );
 a15907a <=( a15906a  and  a15901a );
 a15910a <=( A234  and  A233 );
 a15914a <=( A302  and  A299 );
 a15915a <=( (not A298)  and  a15914a );
 a15916a <=( a15915a  and  a15910a );
 a15919a <=( A166  and  A168 );
 a15923a <=( (not A202)  and  (not A200) );
 a15924a <=( (not A199)  and  a15923a );
 a15925a <=( a15924a  and  a15919a );
 a15928a <=( A234  and  A233 );
 a15932a <=( A269  and  A266 );
 a15933a <=( (not A265)  and  a15932a );
 a15934a <=( a15933a  and  a15928a );
 a15937a <=( A166  and  A168 );
 a15941a <=( (not A202)  and  (not A200) );
 a15942a <=( (not A199)  and  a15941a );
 a15943a <=( a15942a  and  a15937a );
 a15946a <=( A234  and  A233 );
 a15950a <=( A269  and  (not A266) );
 a15951a <=( A265  and  a15950a );
 a15952a <=( a15951a  and  a15946a );
 a15955a <=( A166  and  A168 );
 a15959a <=( (not A202)  and  (not A200) );
 a15960a <=( (not A199)  and  a15959a );
 a15961a <=( a15960a  and  a15955a );
 a15964a <=( A233  and  (not A232) );
 a15968a <=( A300  and  A299 );
 a15969a <=( A236  and  a15968a );
 a15970a <=( a15969a  and  a15964a );
 a15973a <=( A166  and  A168 );
 a15977a <=( (not A202)  and  (not A200) );
 a15978a <=( (not A199)  and  a15977a );
 a15979a <=( a15978a  and  a15973a );
 a15982a <=( A233  and  (not A232) );
 a15986a <=( A300  and  A298 );
 a15987a <=( A236  and  a15986a );
 a15988a <=( a15987a  and  a15982a );
 a15991a <=( A166  and  A168 );
 a15995a <=( (not A202)  and  (not A200) );
 a15996a <=( (not A199)  and  a15995a );
 a15997a <=( a15996a  and  a15991a );
 a16000a <=( A233  and  (not A232) );
 a16004a <=( A267  and  A265 );
 a16005a <=( A236  and  a16004a );
 a16006a <=( a16005a  and  a16000a );
 a16009a <=( A166  and  A168 );
 a16013a <=( (not A202)  and  (not A200) );
 a16014a <=( (not A199)  and  a16013a );
 a16015a <=( a16014a  and  a16009a );
 a16018a <=( A233  and  (not A232) );
 a16022a <=( A267  and  A266 );
 a16023a <=( A236  and  a16022a );
 a16024a <=( a16023a  and  a16018a );
 a16027a <=( A166  and  A168 );
 a16031a <=( (not A202)  and  (not A200) );
 a16032a <=( (not A199)  and  a16031a );
 a16033a <=( a16032a  and  a16027a );
 a16036a <=( (not A233)  and  A232 );
 a16040a <=( A300  and  A299 );
 a16041a <=( A236  and  a16040a );
 a16042a <=( a16041a  and  a16036a );
 a16045a <=( A166  and  A168 );
 a16049a <=( (not A202)  and  (not A200) );
 a16050a <=( (not A199)  and  a16049a );
 a16051a <=( a16050a  and  a16045a );
 a16054a <=( (not A233)  and  A232 );
 a16058a <=( A300  and  A298 );
 a16059a <=( A236  and  a16058a );
 a16060a <=( a16059a  and  a16054a );
 a16063a <=( A166  and  A168 );
 a16067a <=( (not A202)  and  (not A200) );
 a16068a <=( (not A199)  and  a16067a );
 a16069a <=( a16068a  and  a16063a );
 a16072a <=( (not A233)  and  A232 );
 a16076a <=( A267  and  A265 );
 a16077a <=( A236  and  a16076a );
 a16078a <=( a16077a  and  a16072a );
 a16081a <=( A166  and  A168 );
 a16085a <=( (not A202)  and  (not A200) );
 a16086a <=( (not A199)  and  a16085a );
 a16087a <=( a16086a  and  a16081a );
 a16090a <=( (not A233)  and  A232 );
 a16094a <=( A267  and  A266 );
 a16095a <=( A236  and  a16094a );
 a16096a <=( a16095a  and  a16090a );
 a16099a <=( A167  and  A168 );
 a16103a <=( (not A203)  and  (not A202) );
 a16104a <=( (not A201)  and  a16103a );
 a16105a <=( a16104a  and  a16099a );
 a16108a <=( A234  and  A232 );
 a16112a <=( A302  and  (not A299) );
 a16113a <=( A298  and  a16112a );
 a16114a <=( a16113a  and  a16108a );
 a16117a <=( A167  and  A168 );
 a16121a <=( (not A203)  and  (not A202) );
 a16122a <=( (not A201)  and  a16121a );
 a16123a <=( a16122a  and  a16117a );
 a16126a <=( A234  and  A232 );
 a16130a <=( A302  and  A299 );
 a16131a <=( (not A298)  and  a16130a );
 a16132a <=( a16131a  and  a16126a );
 a16135a <=( A167  and  A168 );
 a16139a <=( (not A203)  and  (not A202) );
 a16140a <=( (not A201)  and  a16139a );
 a16141a <=( a16140a  and  a16135a );
 a16144a <=( A234  and  A232 );
 a16148a <=( A269  and  A266 );
 a16149a <=( (not A265)  and  a16148a );
 a16150a <=( a16149a  and  a16144a );
 a16153a <=( A167  and  A168 );
 a16157a <=( (not A203)  and  (not A202) );
 a16158a <=( (not A201)  and  a16157a );
 a16159a <=( a16158a  and  a16153a );
 a16162a <=( A234  and  A232 );
 a16166a <=( A269  and  (not A266) );
 a16167a <=( A265  and  a16166a );
 a16168a <=( a16167a  and  a16162a );
 a16171a <=( A167  and  A168 );
 a16175a <=( (not A203)  and  (not A202) );
 a16176a <=( (not A201)  and  a16175a );
 a16177a <=( a16176a  and  a16171a );
 a16180a <=( A234  and  A233 );
 a16184a <=( A302  and  (not A299) );
 a16185a <=( A298  and  a16184a );
 a16186a <=( a16185a  and  a16180a );
 a16189a <=( A167  and  A168 );
 a16193a <=( (not A203)  and  (not A202) );
 a16194a <=( (not A201)  and  a16193a );
 a16195a <=( a16194a  and  a16189a );
 a16198a <=( A234  and  A233 );
 a16202a <=( A302  and  A299 );
 a16203a <=( (not A298)  and  a16202a );
 a16204a <=( a16203a  and  a16198a );
 a16207a <=( A167  and  A168 );
 a16211a <=( (not A203)  and  (not A202) );
 a16212a <=( (not A201)  and  a16211a );
 a16213a <=( a16212a  and  a16207a );
 a16216a <=( A234  and  A233 );
 a16220a <=( A269  and  A266 );
 a16221a <=( (not A265)  and  a16220a );
 a16222a <=( a16221a  and  a16216a );
 a16225a <=( A167  and  A168 );
 a16229a <=( (not A203)  and  (not A202) );
 a16230a <=( (not A201)  and  a16229a );
 a16231a <=( a16230a  and  a16225a );
 a16234a <=( A234  and  A233 );
 a16238a <=( A269  and  (not A266) );
 a16239a <=( A265  and  a16238a );
 a16240a <=( a16239a  and  a16234a );
 a16243a <=( A167  and  A168 );
 a16247a <=( (not A203)  and  (not A202) );
 a16248a <=( (not A201)  and  a16247a );
 a16249a <=( a16248a  and  a16243a );
 a16252a <=( A233  and  (not A232) );
 a16256a <=( A300  and  A299 );
 a16257a <=( A236  and  a16256a );
 a16258a <=( a16257a  and  a16252a );
 a16261a <=( A167  and  A168 );
 a16265a <=( (not A203)  and  (not A202) );
 a16266a <=( (not A201)  and  a16265a );
 a16267a <=( a16266a  and  a16261a );
 a16270a <=( A233  and  (not A232) );
 a16274a <=( A300  and  A298 );
 a16275a <=( A236  and  a16274a );
 a16276a <=( a16275a  and  a16270a );
 a16279a <=( A167  and  A168 );
 a16283a <=( (not A203)  and  (not A202) );
 a16284a <=( (not A201)  and  a16283a );
 a16285a <=( a16284a  and  a16279a );
 a16288a <=( A233  and  (not A232) );
 a16292a <=( A267  and  A265 );
 a16293a <=( A236  and  a16292a );
 a16294a <=( a16293a  and  a16288a );
 a16297a <=( A167  and  A168 );
 a16301a <=( (not A203)  and  (not A202) );
 a16302a <=( (not A201)  and  a16301a );
 a16303a <=( a16302a  and  a16297a );
 a16306a <=( A233  and  (not A232) );
 a16310a <=( A267  and  A266 );
 a16311a <=( A236  and  a16310a );
 a16312a <=( a16311a  and  a16306a );
 a16315a <=( A167  and  A168 );
 a16319a <=( (not A203)  and  (not A202) );
 a16320a <=( (not A201)  and  a16319a );
 a16321a <=( a16320a  and  a16315a );
 a16324a <=( (not A233)  and  A232 );
 a16328a <=( A300  and  A299 );
 a16329a <=( A236  and  a16328a );
 a16330a <=( a16329a  and  a16324a );
 a16333a <=( A167  and  A168 );
 a16337a <=( (not A203)  and  (not A202) );
 a16338a <=( (not A201)  and  a16337a );
 a16339a <=( a16338a  and  a16333a );
 a16342a <=( (not A233)  and  A232 );
 a16346a <=( A300  and  A298 );
 a16347a <=( A236  and  a16346a );
 a16348a <=( a16347a  and  a16342a );
 a16351a <=( A167  and  A168 );
 a16355a <=( (not A203)  and  (not A202) );
 a16356a <=( (not A201)  and  a16355a );
 a16357a <=( a16356a  and  a16351a );
 a16360a <=( (not A233)  and  A232 );
 a16364a <=( A267  and  A265 );
 a16365a <=( A236  and  a16364a );
 a16366a <=( a16365a  and  a16360a );
 a16369a <=( A167  and  A168 );
 a16373a <=( (not A203)  and  (not A202) );
 a16374a <=( (not A201)  and  a16373a );
 a16375a <=( a16374a  and  a16369a );
 a16378a <=( (not A233)  and  A232 );
 a16382a <=( A267  and  A266 );
 a16383a <=( A236  and  a16382a );
 a16384a <=( a16383a  and  a16378a );
 a16387a <=( A167  and  A168 );
 a16391a <=( (not A201)  and  A200 );
 a16392a <=( A199  and  a16391a );
 a16393a <=( a16392a  and  a16387a );
 a16396a <=( A235  and  (not A202) );
 a16400a <=( A302  and  (not A299) );
 a16401a <=( A298  and  a16400a );
 a16402a <=( a16401a  and  a16396a );
 a16405a <=( A167  and  A168 );
 a16409a <=( (not A201)  and  A200 );
 a16410a <=( A199  and  a16409a );
 a16411a <=( a16410a  and  a16405a );
 a16414a <=( A235  and  (not A202) );
 a16418a <=( A302  and  A299 );
 a16419a <=( (not A298)  and  a16418a );
 a16420a <=( a16419a  and  a16414a );
 a16423a <=( A167  and  A168 );
 a16427a <=( (not A201)  and  A200 );
 a16428a <=( A199  and  a16427a );
 a16429a <=( a16428a  and  a16423a );
 a16432a <=( A235  and  (not A202) );
 a16436a <=( A269  and  A266 );
 a16437a <=( (not A265)  and  a16436a );
 a16438a <=( a16437a  and  a16432a );
 a16441a <=( A167  and  A168 );
 a16445a <=( (not A201)  and  A200 );
 a16446a <=( A199  and  a16445a );
 a16447a <=( a16446a  and  a16441a );
 a16450a <=( A235  and  (not A202) );
 a16454a <=( A269  and  (not A266) );
 a16455a <=( A265  and  a16454a );
 a16456a <=( a16455a  and  a16450a );
 a16459a <=( A167  and  A168 );
 a16463a <=( (not A201)  and  A200 );
 a16464a <=( A199  and  a16463a );
 a16465a <=( a16464a  and  a16459a );
 a16468a <=( A232  and  (not A202) );
 a16472a <=( A300  and  A299 );
 a16473a <=( A234  and  a16472a );
 a16474a <=( a16473a  and  a16468a );
 a16477a <=( A167  and  A168 );
 a16481a <=( (not A201)  and  A200 );
 a16482a <=( A199  and  a16481a );
 a16483a <=( a16482a  and  a16477a );
 a16486a <=( A232  and  (not A202) );
 a16490a <=( A300  and  A298 );
 a16491a <=( A234  and  a16490a );
 a16492a <=( a16491a  and  a16486a );
 a16495a <=( A167  and  A168 );
 a16499a <=( (not A201)  and  A200 );
 a16500a <=( A199  and  a16499a );
 a16501a <=( a16500a  and  a16495a );
 a16504a <=( A232  and  (not A202) );
 a16508a <=( A267  and  A265 );
 a16509a <=( A234  and  a16508a );
 a16510a <=( a16509a  and  a16504a );
 a16513a <=( A167  and  A168 );
 a16517a <=( (not A201)  and  A200 );
 a16518a <=( A199  and  a16517a );
 a16519a <=( a16518a  and  a16513a );
 a16522a <=( A232  and  (not A202) );
 a16526a <=( A267  and  A266 );
 a16527a <=( A234  and  a16526a );
 a16528a <=( a16527a  and  a16522a );
 a16531a <=( A167  and  A168 );
 a16535a <=( (not A201)  and  A200 );
 a16536a <=( A199  and  a16535a );
 a16537a <=( a16536a  and  a16531a );
 a16540a <=( A233  and  (not A202) );
 a16544a <=( A300  and  A299 );
 a16545a <=( A234  and  a16544a );
 a16546a <=( a16545a  and  a16540a );
 a16549a <=( A167  and  A168 );
 a16553a <=( (not A201)  and  A200 );
 a16554a <=( A199  and  a16553a );
 a16555a <=( a16554a  and  a16549a );
 a16558a <=( A233  and  (not A202) );
 a16562a <=( A300  and  A298 );
 a16563a <=( A234  and  a16562a );
 a16564a <=( a16563a  and  a16558a );
 a16567a <=( A167  and  A168 );
 a16571a <=( (not A201)  and  A200 );
 a16572a <=( A199  and  a16571a );
 a16573a <=( a16572a  and  a16567a );
 a16576a <=( A233  and  (not A202) );
 a16580a <=( A267  and  A265 );
 a16581a <=( A234  and  a16580a );
 a16582a <=( a16581a  and  a16576a );
 a16585a <=( A167  and  A168 );
 a16589a <=( (not A201)  and  A200 );
 a16590a <=( A199  and  a16589a );
 a16591a <=( a16590a  and  a16585a );
 a16594a <=( A233  and  (not A202) );
 a16598a <=( A267  and  A266 );
 a16599a <=( A234  and  a16598a );
 a16600a <=( a16599a  and  a16594a );
 a16603a <=( A167  and  A168 );
 a16607a <=( (not A201)  and  A200 );
 a16608a <=( A199  and  a16607a );
 a16609a <=( a16608a  and  a16603a );
 a16612a <=( (not A232)  and  (not A202) );
 a16616a <=( A301  and  A236 );
 a16617a <=( A233  and  a16616a );
 a16618a <=( a16617a  and  a16612a );
 a16621a <=( A167  and  A168 );
 a16625a <=( (not A201)  and  A200 );
 a16626a <=( A199  and  a16625a );
 a16627a <=( a16626a  and  a16621a );
 a16630a <=( (not A232)  and  (not A202) );
 a16634a <=( A268  and  A236 );
 a16635a <=( A233  and  a16634a );
 a16636a <=( a16635a  and  a16630a );
 a16639a <=( A167  and  A168 );
 a16643a <=( (not A201)  and  A200 );
 a16644a <=( A199  and  a16643a );
 a16645a <=( a16644a  and  a16639a );
 a16648a <=( A232  and  (not A202) );
 a16652a <=( A301  and  A236 );
 a16653a <=( (not A233)  and  a16652a );
 a16654a <=( a16653a  and  a16648a );
 a16657a <=( A167  and  A168 );
 a16661a <=( (not A201)  and  A200 );
 a16662a <=( A199  and  a16661a );
 a16663a <=( a16662a  and  a16657a );
 a16666a <=( A232  and  (not A202) );
 a16670a <=( A268  and  A236 );
 a16671a <=( (not A233)  and  a16670a );
 a16672a <=( a16671a  and  a16666a );
 a16675a <=( A167  and  A168 );
 a16679a <=( (not A202)  and  (not A200) );
 a16680a <=( (not A199)  and  a16679a );
 a16681a <=( a16680a  and  a16675a );
 a16684a <=( A234  and  A232 );
 a16688a <=( A302  and  (not A299) );
 a16689a <=( A298  and  a16688a );
 a16690a <=( a16689a  and  a16684a );
 a16693a <=( A167  and  A168 );
 a16697a <=( (not A202)  and  (not A200) );
 a16698a <=( (not A199)  and  a16697a );
 a16699a <=( a16698a  and  a16693a );
 a16702a <=( A234  and  A232 );
 a16706a <=( A302  and  A299 );
 a16707a <=( (not A298)  and  a16706a );
 a16708a <=( a16707a  and  a16702a );
 a16711a <=( A167  and  A168 );
 a16715a <=( (not A202)  and  (not A200) );
 a16716a <=( (not A199)  and  a16715a );
 a16717a <=( a16716a  and  a16711a );
 a16720a <=( A234  and  A232 );
 a16724a <=( A269  and  A266 );
 a16725a <=( (not A265)  and  a16724a );
 a16726a <=( a16725a  and  a16720a );
 a16729a <=( A167  and  A168 );
 a16733a <=( (not A202)  and  (not A200) );
 a16734a <=( (not A199)  and  a16733a );
 a16735a <=( a16734a  and  a16729a );
 a16738a <=( A234  and  A232 );
 a16742a <=( A269  and  (not A266) );
 a16743a <=( A265  and  a16742a );
 a16744a <=( a16743a  and  a16738a );
 a16747a <=( A167  and  A168 );
 a16751a <=( (not A202)  and  (not A200) );
 a16752a <=( (not A199)  and  a16751a );
 a16753a <=( a16752a  and  a16747a );
 a16756a <=( A234  and  A233 );
 a16760a <=( A302  and  (not A299) );
 a16761a <=( A298  and  a16760a );
 a16762a <=( a16761a  and  a16756a );
 a16765a <=( A167  and  A168 );
 a16769a <=( (not A202)  and  (not A200) );
 a16770a <=( (not A199)  and  a16769a );
 a16771a <=( a16770a  and  a16765a );
 a16774a <=( A234  and  A233 );
 a16778a <=( A302  and  A299 );
 a16779a <=( (not A298)  and  a16778a );
 a16780a <=( a16779a  and  a16774a );
 a16783a <=( A167  and  A168 );
 a16787a <=( (not A202)  and  (not A200) );
 a16788a <=( (not A199)  and  a16787a );
 a16789a <=( a16788a  and  a16783a );
 a16792a <=( A234  and  A233 );
 a16796a <=( A269  and  A266 );
 a16797a <=( (not A265)  and  a16796a );
 a16798a <=( a16797a  and  a16792a );
 a16801a <=( A167  and  A168 );
 a16805a <=( (not A202)  and  (not A200) );
 a16806a <=( (not A199)  and  a16805a );
 a16807a <=( a16806a  and  a16801a );
 a16810a <=( A234  and  A233 );
 a16814a <=( A269  and  (not A266) );
 a16815a <=( A265  and  a16814a );
 a16816a <=( a16815a  and  a16810a );
 a16819a <=( A167  and  A168 );
 a16823a <=( (not A202)  and  (not A200) );
 a16824a <=( (not A199)  and  a16823a );
 a16825a <=( a16824a  and  a16819a );
 a16828a <=( A233  and  (not A232) );
 a16832a <=( A300  and  A299 );
 a16833a <=( A236  and  a16832a );
 a16834a <=( a16833a  and  a16828a );
 a16837a <=( A167  and  A168 );
 a16841a <=( (not A202)  and  (not A200) );
 a16842a <=( (not A199)  and  a16841a );
 a16843a <=( a16842a  and  a16837a );
 a16846a <=( A233  and  (not A232) );
 a16850a <=( A300  and  A298 );
 a16851a <=( A236  and  a16850a );
 a16852a <=( a16851a  and  a16846a );
 a16855a <=( A167  and  A168 );
 a16859a <=( (not A202)  and  (not A200) );
 a16860a <=( (not A199)  and  a16859a );
 a16861a <=( a16860a  and  a16855a );
 a16864a <=( A233  and  (not A232) );
 a16868a <=( A267  and  A265 );
 a16869a <=( A236  and  a16868a );
 a16870a <=( a16869a  and  a16864a );
 a16873a <=( A167  and  A168 );
 a16877a <=( (not A202)  and  (not A200) );
 a16878a <=( (not A199)  and  a16877a );
 a16879a <=( a16878a  and  a16873a );
 a16882a <=( A233  and  (not A232) );
 a16886a <=( A267  and  A266 );
 a16887a <=( A236  and  a16886a );
 a16888a <=( a16887a  and  a16882a );
 a16891a <=( A167  and  A168 );
 a16895a <=( (not A202)  and  (not A200) );
 a16896a <=( (not A199)  and  a16895a );
 a16897a <=( a16896a  and  a16891a );
 a16900a <=( (not A233)  and  A232 );
 a16904a <=( A300  and  A299 );
 a16905a <=( A236  and  a16904a );
 a16906a <=( a16905a  and  a16900a );
 a16909a <=( A167  and  A168 );
 a16913a <=( (not A202)  and  (not A200) );
 a16914a <=( (not A199)  and  a16913a );
 a16915a <=( a16914a  and  a16909a );
 a16918a <=( (not A233)  and  A232 );
 a16922a <=( A300  and  A298 );
 a16923a <=( A236  and  a16922a );
 a16924a <=( a16923a  and  a16918a );
 a16927a <=( A167  and  A168 );
 a16931a <=( (not A202)  and  (not A200) );
 a16932a <=( (not A199)  and  a16931a );
 a16933a <=( a16932a  and  a16927a );
 a16936a <=( (not A233)  and  A232 );
 a16940a <=( A267  and  A265 );
 a16941a <=( A236  and  a16940a );
 a16942a <=( a16941a  and  a16936a );
 a16945a <=( A167  and  A168 );
 a16949a <=( (not A202)  and  (not A200) );
 a16950a <=( (not A199)  and  a16949a );
 a16951a <=( a16950a  and  a16945a );
 a16954a <=( (not A233)  and  A232 );
 a16958a <=( A267  and  A266 );
 a16959a <=( A236  and  a16958a );
 a16960a <=( a16959a  and  a16954a );
 a16963a <=( A167  and  A170 );
 a16967a <=( (not A202)  and  (not A201) );
 a16968a <=( (not A166)  and  a16967a );
 a16969a <=( a16968a  and  a16963a );
 a16972a <=( A235  and  (not A203) );
 a16976a <=( A302  and  (not A299) );
 a16977a <=( A298  and  a16976a );
 a16978a <=( a16977a  and  a16972a );
 a16981a <=( A167  and  A170 );
 a16985a <=( (not A202)  and  (not A201) );
 a16986a <=( (not A166)  and  a16985a );
 a16987a <=( a16986a  and  a16981a );
 a16990a <=( A235  and  (not A203) );
 a16994a <=( A302  and  A299 );
 a16995a <=( (not A298)  and  a16994a );
 a16996a <=( a16995a  and  a16990a );
 a16999a <=( A167  and  A170 );
 a17003a <=( (not A202)  and  (not A201) );
 a17004a <=( (not A166)  and  a17003a );
 a17005a <=( a17004a  and  a16999a );
 a17008a <=( A235  and  (not A203) );
 a17012a <=( A269  and  A266 );
 a17013a <=( (not A265)  and  a17012a );
 a17014a <=( a17013a  and  a17008a );
 a17017a <=( A167  and  A170 );
 a17021a <=( (not A202)  and  (not A201) );
 a17022a <=( (not A166)  and  a17021a );
 a17023a <=( a17022a  and  a17017a );
 a17026a <=( A235  and  (not A203) );
 a17030a <=( A269  and  (not A266) );
 a17031a <=( A265  and  a17030a );
 a17032a <=( a17031a  and  a17026a );
 a17035a <=( A167  and  A170 );
 a17039a <=( (not A202)  and  (not A201) );
 a17040a <=( (not A166)  and  a17039a );
 a17041a <=( a17040a  and  a17035a );
 a17044a <=( A232  and  (not A203) );
 a17048a <=( A300  and  A299 );
 a17049a <=( A234  and  a17048a );
 a17050a <=( a17049a  and  a17044a );
 a17053a <=( A167  and  A170 );
 a17057a <=( (not A202)  and  (not A201) );
 a17058a <=( (not A166)  and  a17057a );
 a17059a <=( a17058a  and  a17053a );
 a17062a <=( A232  and  (not A203) );
 a17066a <=( A300  and  A298 );
 a17067a <=( A234  and  a17066a );
 a17068a <=( a17067a  and  a17062a );
 a17071a <=( A167  and  A170 );
 a17075a <=( (not A202)  and  (not A201) );
 a17076a <=( (not A166)  and  a17075a );
 a17077a <=( a17076a  and  a17071a );
 a17080a <=( A232  and  (not A203) );
 a17084a <=( A267  and  A265 );
 a17085a <=( A234  and  a17084a );
 a17086a <=( a17085a  and  a17080a );
 a17089a <=( A167  and  A170 );
 a17093a <=( (not A202)  and  (not A201) );
 a17094a <=( (not A166)  and  a17093a );
 a17095a <=( a17094a  and  a17089a );
 a17098a <=( A232  and  (not A203) );
 a17102a <=( A267  and  A266 );
 a17103a <=( A234  and  a17102a );
 a17104a <=( a17103a  and  a17098a );
 a17107a <=( A167  and  A170 );
 a17111a <=( (not A202)  and  (not A201) );
 a17112a <=( (not A166)  and  a17111a );
 a17113a <=( a17112a  and  a17107a );
 a17116a <=( A233  and  (not A203) );
 a17120a <=( A300  and  A299 );
 a17121a <=( A234  and  a17120a );
 a17122a <=( a17121a  and  a17116a );
 a17125a <=( A167  and  A170 );
 a17129a <=( (not A202)  and  (not A201) );
 a17130a <=( (not A166)  and  a17129a );
 a17131a <=( a17130a  and  a17125a );
 a17134a <=( A233  and  (not A203) );
 a17138a <=( A300  and  A298 );
 a17139a <=( A234  and  a17138a );
 a17140a <=( a17139a  and  a17134a );
 a17143a <=( A167  and  A170 );
 a17147a <=( (not A202)  and  (not A201) );
 a17148a <=( (not A166)  and  a17147a );
 a17149a <=( a17148a  and  a17143a );
 a17152a <=( A233  and  (not A203) );
 a17156a <=( A267  and  A265 );
 a17157a <=( A234  and  a17156a );
 a17158a <=( a17157a  and  a17152a );
 a17161a <=( A167  and  A170 );
 a17165a <=( (not A202)  and  (not A201) );
 a17166a <=( (not A166)  and  a17165a );
 a17167a <=( a17166a  and  a17161a );
 a17170a <=( A233  and  (not A203) );
 a17174a <=( A267  and  A266 );
 a17175a <=( A234  and  a17174a );
 a17176a <=( a17175a  and  a17170a );
 a17179a <=( A167  and  A170 );
 a17183a <=( (not A202)  and  (not A201) );
 a17184a <=( (not A166)  and  a17183a );
 a17185a <=( a17184a  and  a17179a );
 a17188a <=( (not A232)  and  (not A203) );
 a17192a <=( A301  and  A236 );
 a17193a <=( A233  and  a17192a );
 a17194a <=( a17193a  and  a17188a );
 a17197a <=( A167  and  A170 );
 a17201a <=( (not A202)  and  (not A201) );
 a17202a <=( (not A166)  and  a17201a );
 a17203a <=( a17202a  and  a17197a );
 a17206a <=( (not A232)  and  (not A203) );
 a17210a <=( A268  and  A236 );
 a17211a <=( A233  and  a17210a );
 a17212a <=( a17211a  and  a17206a );
 a17215a <=( A167  and  A170 );
 a17219a <=( (not A202)  and  (not A201) );
 a17220a <=( (not A166)  and  a17219a );
 a17221a <=( a17220a  and  a17215a );
 a17224a <=( A232  and  (not A203) );
 a17228a <=( A301  and  A236 );
 a17229a <=( (not A233)  and  a17228a );
 a17230a <=( a17229a  and  a17224a );
 a17233a <=( A167  and  A170 );
 a17237a <=( (not A202)  and  (not A201) );
 a17238a <=( (not A166)  and  a17237a );
 a17239a <=( a17238a  and  a17233a );
 a17242a <=( A232  and  (not A203) );
 a17246a <=( A268  and  A236 );
 a17247a <=( (not A233)  and  a17246a );
 a17248a <=( a17247a  and  a17242a );
 a17251a <=( A167  and  A170 );
 a17255a <=( A200  and  A199 );
 a17256a <=( (not A166)  and  a17255a );
 a17257a <=( a17256a  and  a17251a );
 a17260a <=( (not A202)  and  (not A201) );
 a17264a <=( A300  and  A299 );
 a17265a <=( A235  and  a17264a );
 a17266a <=( a17265a  and  a17260a );
 a17269a <=( A167  and  A170 );
 a17273a <=( A200  and  A199 );
 a17274a <=( (not A166)  and  a17273a );
 a17275a <=( a17274a  and  a17269a );
 a17278a <=( (not A202)  and  (not A201) );
 a17282a <=( A300  and  A298 );
 a17283a <=( A235  and  a17282a );
 a17284a <=( a17283a  and  a17278a );
 a17287a <=( A167  and  A170 );
 a17291a <=( A200  and  A199 );
 a17292a <=( (not A166)  and  a17291a );
 a17293a <=( a17292a  and  a17287a );
 a17296a <=( (not A202)  and  (not A201) );
 a17300a <=( A267  and  A265 );
 a17301a <=( A235  and  a17300a );
 a17302a <=( a17301a  and  a17296a );
 a17305a <=( A167  and  A170 );
 a17309a <=( A200  and  A199 );
 a17310a <=( (not A166)  and  a17309a );
 a17311a <=( a17310a  and  a17305a );
 a17314a <=( (not A202)  and  (not A201) );
 a17318a <=( A267  and  A266 );
 a17319a <=( A235  and  a17318a );
 a17320a <=( a17319a  and  a17314a );
 a17323a <=( A167  and  A170 );
 a17327a <=( A200  and  A199 );
 a17328a <=( (not A166)  and  a17327a );
 a17329a <=( a17328a  and  a17323a );
 a17332a <=( (not A202)  and  (not A201) );
 a17336a <=( A301  and  A234 );
 a17337a <=( A232  and  a17336a );
 a17338a <=( a17337a  and  a17332a );
 a17341a <=( A167  and  A170 );
 a17345a <=( A200  and  A199 );
 a17346a <=( (not A166)  and  a17345a );
 a17347a <=( a17346a  and  a17341a );
 a17350a <=( (not A202)  and  (not A201) );
 a17354a <=( A268  and  A234 );
 a17355a <=( A232  and  a17354a );
 a17356a <=( a17355a  and  a17350a );
 a17359a <=( A167  and  A170 );
 a17363a <=( A200  and  A199 );
 a17364a <=( (not A166)  and  a17363a );
 a17365a <=( a17364a  and  a17359a );
 a17368a <=( (not A202)  and  (not A201) );
 a17372a <=( A301  and  A234 );
 a17373a <=( A233  and  a17372a );
 a17374a <=( a17373a  and  a17368a );
 a17377a <=( A167  and  A170 );
 a17381a <=( A200  and  A199 );
 a17382a <=( (not A166)  and  a17381a );
 a17383a <=( a17382a  and  a17377a );
 a17386a <=( (not A202)  and  (not A201) );
 a17390a <=( A268  and  A234 );
 a17391a <=( A233  and  a17390a );
 a17392a <=( a17391a  and  a17386a );
 a17395a <=( A167  and  A170 );
 a17399a <=( (not A200)  and  (not A199) );
 a17400a <=( (not A166)  and  a17399a );
 a17401a <=( a17400a  and  a17395a );
 a17404a <=( A235  and  (not A202) );
 a17408a <=( A302  and  (not A299) );
 a17409a <=( A298  and  a17408a );
 a17410a <=( a17409a  and  a17404a );
 a17413a <=( A167  and  A170 );
 a17417a <=( (not A200)  and  (not A199) );
 a17418a <=( (not A166)  and  a17417a );
 a17419a <=( a17418a  and  a17413a );
 a17422a <=( A235  and  (not A202) );
 a17426a <=( A302  and  A299 );
 a17427a <=( (not A298)  and  a17426a );
 a17428a <=( a17427a  and  a17422a );
 a17431a <=( A167  and  A170 );
 a17435a <=( (not A200)  and  (not A199) );
 a17436a <=( (not A166)  and  a17435a );
 a17437a <=( a17436a  and  a17431a );
 a17440a <=( A235  and  (not A202) );
 a17444a <=( A269  and  A266 );
 a17445a <=( (not A265)  and  a17444a );
 a17446a <=( a17445a  and  a17440a );
 a17449a <=( A167  and  A170 );
 a17453a <=( (not A200)  and  (not A199) );
 a17454a <=( (not A166)  and  a17453a );
 a17455a <=( a17454a  and  a17449a );
 a17458a <=( A235  and  (not A202) );
 a17462a <=( A269  and  (not A266) );
 a17463a <=( A265  and  a17462a );
 a17464a <=( a17463a  and  a17458a );
 a17467a <=( A167  and  A170 );
 a17471a <=( (not A200)  and  (not A199) );
 a17472a <=( (not A166)  and  a17471a );
 a17473a <=( a17472a  and  a17467a );
 a17476a <=( A232  and  (not A202) );
 a17480a <=( A300  and  A299 );
 a17481a <=( A234  and  a17480a );
 a17482a <=( a17481a  and  a17476a );
 a17485a <=( A167  and  A170 );
 a17489a <=( (not A200)  and  (not A199) );
 a17490a <=( (not A166)  and  a17489a );
 a17491a <=( a17490a  and  a17485a );
 a17494a <=( A232  and  (not A202) );
 a17498a <=( A300  and  A298 );
 a17499a <=( A234  and  a17498a );
 a17500a <=( a17499a  and  a17494a );
 a17503a <=( A167  and  A170 );
 a17507a <=( (not A200)  and  (not A199) );
 a17508a <=( (not A166)  and  a17507a );
 a17509a <=( a17508a  and  a17503a );
 a17512a <=( A232  and  (not A202) );
 a17516a <=( A267  and  A265 );
 a17517a <=( A234  and  a17516a );
 a17518a <=( a17517a  and  a17512a );
 a17521a <=( A167  and  A170 );
 a17525a <=( (not A200)  and  (not A199) );
 a17526a <=( (not A166)  and  a17525a );
 a17527a <=( a17526a  and  a17521a );
 a17530a <=( A232  and  (not A202) );
 a17534a <=( A267  and  A266 );
 a17535a <=( A234  and  a17534a );
 a17536a <=( a17535a  and  a17530a );
 a17539a <=( A167  and  A170 );
 a17543a <=( (not A200)  and  (not A199) );
 a17544a <=( (not A166)  and  a17543a );
 a17545a <=( a17544a  and  a17539a );
 a17548a <=( A233  and  (not A202) );
 a17552a <=( A300  and  A299 );
 a17553a <=( A234  and  a17552a );
 a17554a <=( a17553a  and  a17548a );
 a17557a <=( A167  and  A170 );
 a17561a <=( (not A200)  and  (not A199) );
 a17562a <=( (not A166)  and  a17561a );
 a17563a <=( a17562a  and  a17557a );
 a17566a <=( A233  and  (not A202) );
 a17570a <=( A300  and  A298 );
 a17571a <=( A234  and  a17570a );
 a17572a <=( a17571a  and  a17566a );
 a17575a <=( A167  and  A170 );
 a17579a <=( (not A200)  and  (not A199) );
 a17580a <=( (not A166)  and  a17579a );
 a17581a <=( a17580a  and  a17575a );
 a17584a <=( A233  and  (not A202) );
 a17588a <=( A267  and  A265 );
 a17589a <=( A234  and  a17588a );
 a17590a <=( a17589a  and  a17584a );
 a17593a <=( A167  and  A170 );
 a17597a <=( (not A200)  and  (not A199) );
 a17598a <=( (not A166)  and  a17597a );
 a17599a <=( a17598a  and  a17593a );
 a17602a <=( A233  and  (not A202) );
 a17606a <=( A267  and  A266 );
 a17607a <=( A234  and  a17606a );
 a17608a <=( a17607a  and  a17602a );
 a17611a <=( A167  and  A170 );
 a17615a <=( (not A200)  and  (not A199) );
 a17616a <=( (not A166)  and  a17615a );
 a17617a <=( a17616a  and  a17611a );
 a17620a <=( (not A232)  and  (not A202) );
 a17624a <=( A301  and  A236 );
 a17625a <=( A233  and  a17624a );
 a17626a <=( a17625a  and  a17620a );
 a17629a <=( A167  and  A170 );
 a17633a <=( (not A200)  and  (not A199) );
 a17634a <=( (not A166)  and  a17633a );
 a17635a <=( a17634a  and  a17629a );
 a17638a <=( (not A232)  and  (not A202) );
 a17642a <=( A268  and  A236 );
 a17643a <=( A233  and  a17642a );
 a17644a <=( a17643a  and  a17638a );
 a17647a <=( A167  and  A170 );
 a17651a <=( (not A200)  and  (not A199) );
 a17652a <=( (not A166)  and  a17651a );
 a17653a <=( a17652a  and  a17647a );
 a17656a <=( A232  and  (not A202) );
 a17660a <=( A301  and  A236 );
 a17661a <=( (not A233)  and  a17660a );
 a17662a <=( a17661a  and  a17656a );
 a17665a <=( A167  and  A170 );
 a17669a <=( (not A200)  and  (not A199) );
 a17670a <=( (not A166)  and  a17669a );
 a17671a <=( a17670a  and  a17665a );
 a17674a <=( A232  and  (not A202) );
 a17678a <=( A268  and  A236 );
 a17679a <=( (not A233)  and  a17678a );
 a17680a <=( a17679a  and  a17674a );
 a17683a <=( (not A167)  and  A170 );
 a17687a <=( (not A202)  and  (not A201) );
 a17688a <=( A166  and  a17687a );
 a17689a <=( a17688a  and  a17683a );
 a17692a <=( A235  and  (not A203) );
 a17696a <=( A302  and  (not A299) );
 a17697a <=( A298  and  a17696a );
 a17698a <=( a17697a  and  a17692a );
 a17701a <=( (not A167)  and  A170 );
 a17705a <=( (not A202)  and  (not A201) );
 a17706a <=( A166  and  a17705a );
 a17707a <=( a17706a  and  a17701a );
 a17710a <=( A235  and  (not A203) );
 a17714a <=( A302  and  A299 );
 a17715a <=( (not A298)  and  a17714a );
 a17716a <=( a17715a  and  a17710a );
 a17719a <=( (not A167)  and  A170 );
 a17723a <=( (not A202)  and  (not A201) );
 a17724a <=( A166  and  a17723a );
 a17725a <=( a17724a  and  a17719a );
 a17728a <=( A235  and  (not A203) );
 a17732a <=( A269  and  A266 );
 a17733a <=( (not A265)  and  a17732a );
 a17734a <=( a17733a  and  a17728a );
 a17737a <=( (not A167)  and  A170 );
 a17741a <=( (not A202)  and  (not A201) );
 a17742a <=( A166  and  a17741a );
 a17743a <=( a17742a  and  a17737a );
 a17746a <=( A235  and  (not A203) );
 a17750a <=( A269  and  (not A266) );
 a17751a <=( A265  and  a17750a );
 a17752a <=( a17751a  and  a17746a );
 a17755a <=( (not A167)  and  A170 );
 a17759a <=( (not A202)  and  (not A201) );
 a17760a <=( A166  and  a17759a );
 a17761a <=( a17760a  and  a17755a );
 a17764a <=( A232  and  (not A203) );
 a17768a <=( A300  and  A299 );
 a17769a <=( A234  and  a17768a );
 a17770a <=( a17769a  and  a17764a );
 a17773a <=( (not A167)  and  A170 );
 a17777a <=( (not A202)  and  (not A201) );
 a17778a <=( A166  and  a17777a );
 a17779a <=( a17778a  and  a17773a );
 a17782a <=( A232  and  (not A203) );
 a17786a <=( A300  and  A298 );
 a17787a <=( A234  and  a17786a );
 a17788a <=( a17787a  and  a17782a );
 a17791a <=( (not A167)  and  A170 );
 a17795a <=( (not A202)  and  (not A201) );
 a17796a <=( A166  and  a17795a );
 a17797a <=( a17796a  and  a17791a );
 a17800a <=( A232  and  (not A203) );
 a17804a <=( A267  and  A265 );
 a17805a <=( A234  and  a17804a );
 a17806a <=( a17805a  and  a17800a );
 a17809a <=( (not A167)  and  A170 );
 a17813a <=( (not A202)  and  (not A201) );
 a17814a <=( A166  and  a17813a );
 a17815a <=( a17814a  and  a17809a );
 a17818a <=( A232  and  (not A203) );
 a17822a <=( A267  and  A266 );
 a17823a <=( A234  and  a17822a );
 a17824a <=( a17823a  and  a17818a );
 a17827a <=( (not A167)  and  A170 );
 a17831a <=( (not A202)  and  (not A201) );
 a17832a <=( A166  and  a17831a );
 a17833a <=( a17832a  and  a17827a );
 a17836a <=( A233  and  (not A203) );
 a17840a <=( A300  and  A299 );
 a17841a <=( A234  and  a17840a );
 a17842a <=( a17841a  and  a17836a );
 a17845a <=( (not A167)  and  A170 );
 a17849a <=( (not A202)  and  (not A201) );
 a17850a <=( A166  and  a17849a );
 a17851a <=( a17850a  and  a17845a );
 a17854a <=( A233  and  (not A203) );
 a17858a <=( A300  and  A298 );
 a17859a <=( A234  and  a17858a );
 a17860a <=( a17859a  and  a17854a );
 a17863a <=( (not A167)  and  A170 );
 a17867a <=( (not A202)  and  (not A201) );
 a17868a <=( A166  and  a17867a );
 a17869a <=( a17868a  and  a17863a );
 a17872a <=( A233  and  (not A203) );
 a17876a <=( A267  and  A265 );
 a17877a <=( A234  and  a17876a );
 a17878a <=( a17877a  and  a17872a );
 a17881a <=( (not A167)  and  A170 );
 a17885a <=( (not A202)  and  (not A201) );
 a17886a <=( A166  and  a17885a );
 a17887a <=( a17886a  and  a17881a );
 a17890a <=( A233  and  (not A203) );
 a17894a <=( A267  and  A266 );
 a17895a <=( A234  and  a17894a );
 a17896a <=( a17895a  and  a17890a );
 a17899a <=( (not A167)  and  A170 );
 a17903a <=( (not A202)  and  (not A201) );
 a17904a <=( A166  and  a17903a );
 a17905a <=( a17904a  and  a17899a );
 a17908a <=( (not A232)  and  (not A203) );
 a17912a <=( A301  and  A236 );
 a17913a <=( A233  and  a17912a );
 a17914a <=( a17913a  and  a17908a );
 a17917a <=( (not A167)  and  A170 );
 a17921a <=( (not A202)  and  (not A201) );
 a17922a <=( A166  and  a17921a );
 a17923a <=( a17922a  and  a17917a );
 a17926a <=( (not A232)  and  (not A203) );
 a17930a <=( A268  and  A236 );
 a17931a <=( A233  and  a17930a );
 a17932a <=( a17931a  and  a17926a );
 a17935a <=( (not A167)  and  A170 );
 a17939a <=( (not A202)  and  (not A201) );
 a17940a <=( A166  and  a17939a );
 a17941a <=( a17940a  and  a17935a );
 a17944a <=( A232  and  (not A203) );
 a17948a <=( A301  and  A236 );
 a17949a <=( (not A233)  and  a17948a );
 a17950a <=( a17949a  and  a17944a );
 a17953a <=( (not A167)  and  A170 );
 a17957a <=( (not A202)  and  (not A201) );
 a17958a <=( A166  and  a17957a );
 a17959a <=( a17958a  and  a17953a );
 a17962a <=( A232  and  (not A203) );
 a17966a <=( A268  and  A236 );
 a17967a <=( (not A233)  and  a17966a );
 a17968a <=( a17967a  and  a17962a );
 a17971a <=( (not A167)  and  A170 );
 a17975a <=( A200  and  A199 );
 a17976a <=( A166  and  a17975a );
 a17977a <=( a17976a  and  a17971a );
 a17980a <=( (not A202)  and  (not A201) );
 a17984a <=( A300  and  A299 );
 a17985a <=( A235  and  a17984a );
 a17986a <=( a17985a  and  a17980a );
 a17989a <=( (not A167)  and  A170 );
 a17993a <=( A200  and  A199 );
 a17994a <=( A166  and  a17993a );
 a17995a <=( a17994a  and  a17989a );
 a17998a <=( (not A202)  and  (not A201) );
 a18002a <=( A300  and  A298 );
 a18003a <=( A235  and  a18002a );
 a18004a <=( a18003a  and  a17998a );
 a18007a <=( (not A167)  and  A170 );
 a18011a <=( A200  and  A199 );
 a18012a <=( A166  and  a18011a );
 a18013a <=( a18012a  and  a18007a );
 a18016a <=( (not A202)  and  (not A201) );
 a18020a <=( A267  and  A265 );
 a18021a <=( A235  and  a18020a );
 a18022a <=( a18021a  and  a18016a );
 a18025a <=( (not A167)  and  A170 );
 a18029a <=( A200  and  A199 );
 a18030a <=( A166  and  a18029a );
 a18031a <=( a18030a  and  a18025a );
 a18034a <=( (not A202)  and  (not A201) );
 a18038a <=( A267  and  A266 );
 a18039a <=( A235  and  a18038a );
 a18040a <=( a18039a  and  a18034a );
 a18043a <=( (not A167)  and  A170 );
 a18047a <=( A200  and  A199 );
 a18048a <=( A166  and  a18047a );
 a18049a <=( a18048a  and  a18043a );
 a18052a <=( (not A202)  and  (not A201) );
 a18056a <=( A301  and  A234 );
 a18057a <=( A232  and  a18056a );
 a18058a <=( a18057a  and  a18052a );
 a18061a <=( (not A167)  and  A170 );
 a18065a <=( A200  and  A199 );
 a18066a <=( A166  and  a18065a );
 a18067a <=( a18066a  and  a18061a );
 a18070a <=( (not A202)  and  (not A201) );
 a18074a <=( A268  and  A234 );
 a18075a <=( A232  and  a18074a );
 a18076a <=( a18075a  and  a18070a );
 a18079a <=( (not A167)  and  A170 );
 a18083a <=( A200  and  A199 );
 a18084a <=( A166  and  a18083a );
 a18085a <=( a18084a  and  a18079a );
 a18088a <=( (not A202)  and  (not A201) );
 a18092a <=( A301  and  A234 );
 a18093a <=( A233  and  a18092a );
 a18094a <=( a18093a  and  a18088a );
 a18097a <=( (not A167)  and  A170 );
 a18101a <=( A200  and  A199 );
 a18102a <=( A166  and  a18101a );
 a18103a <=( a18102a  and  a18097a );
 a18106a <=( (not A202)  and  (not A201) );
 a18110a <=( A268  and  A234 );
 a18111a <=( A233  and  a18110a );
 a18112a <=( a18111a  and  a18106a );
 a18115a <=( (not A167)  and  A170 );
 a18119a <=( (not A200)  and  (not A199) );
 a18120a <=( A166  and  a18119a );
 a18121a <=( a18120a  and  a18115a );
 a18124a <=( A235  and  (not A202) );
 a18128a <=( A302  and  (not A299) );
 a18129a <=( A298  and  a18128a );
 a18130a <=( a18129a  and  a18124a );
 a18133a <=( (not A167)  and  A170 );
 a18137a <=( (not A200)  and  (not A199) );
 a18138a <=( A166  and  a18137a );
 a18139a <=( a18138a  and  a18133a );
 a18142a <=( A235  and  (not A202) );
 a18146a <=( A302  and  A299 );
 a18147a <=( (not A298)  and  a18146a );
 a18148a <=( a18147a  and  a18142a );
 a18151a <=( (not A167)  and  A170 );
 a18155a <=( (not A200)  and  (not A199) );
 a18156a <=( A166  and  a18155a );
 a18157a <=( a18156a  and  a18151a );
 a18160a <=( A235  and  (not A202) );
 a18164a <=( A269  and  A266 );
 a18165a <=( (not A265)  and  a18164a );
 a18166a <=( a18165a  and  a18160a );
 a18169a <=( (not A167)  and  A170 );
 a18173a <=( (not A200)  and  (not A199) );
 a18174a <=( A166  and  a18173a );
 a18175a <=( a18174a  and  a18169a );
 a18178a <=( A235  and  (not A202) );
 a18182a <=( A269  and  (not A266) );
 a18183a <=( A265  and  a18182a );
 a18184a <=( a18183a  and  a18178a );
 a18187a <=( (not A167)  and  A170 );
 a18191a <=( (not A200)  and  (not A199) );
 a18192a <=( A166  and  a18191a );
 a18193a <=( a18192a  and  a18187a );
 a18196a <=( A232  and  (not A202) );
 a18200a <=( A300  and  A299 );
 a18201a <=( A234  and  a18200a );
 a18202a <=( a18201a  and  a18196a );
 a18205a <=( (not A167)  and  A170 );
 a18209a <=( (not A200)  and  (not A199) );
 a18210a <=( A166  and  a18209a );
 a18211a <=( a18210a  and  a18205a );
 a18214a <=( A232  and  (not A202) );
 a18218a <=( A300  and  A298 );
 a18219a <=( A234  and  a18218a );
 a18220a <=( a18219a  and  a18214a );
 a18223a <=( (not A167)  and  A170 );
 a18227a <=( (not A200)  and  (not A199) );
 a18228a <=( A166  and  a18227a );
 a18229a <=( a18228a  and  a18223a );
 a18232a <=( A232  and  (not A202) );
 a18236a <=( A267  and  A265 );
 a18237a <=( A234  and  a18236a );
 a18238a <=( a18237a  and  a18232a );
 a18241a <=( (not A167)  and  A170 );
 a18245a <=( (not A200)  and  (not A199) );
 a18246a <=( A166  and  a18245a );
 a18247a <=( a18246a  and  a18241a );
 a18250a <=( A232  and  (not A202) );
 a18254a <=( A267  and  A266 );
 a18255a <=( A234  and  a18254a );
 a18256a <=( a18255a  and  a18250a );
 a18259a <=( (not A167)  and  A170 );
 a18263a <=( (not A200)  and  (not A199) );
 a18264a <=( A166  and  a18263a );
 a18265a <=( a18264a  and  a18259a );
 a18268a <=( A233  and  (not A202) );
 a18272a <=( A300  and  A299 );
 a18273a <=( A234  and  a18272a );
 a18274a <=( a18273a  and  a18268a );
 a18277a <=( (not A167)  and  A170 );
 a18281a <=( (not A200)  and  (not A199) );
 a18282a <=( A166  and  a18281a );
 a18283a <=( a18282a  and  a18277a );
 a18286a <=( A233  and  (not A202) );
 a18290a <=( A300  and  A298 );
 a18291a <=( A234  and  a18290a );
 a18292a <=( a18291a  and  a18286a );
 a18295a <=( (not A167)  and  A170 );
 a18299a <=( (not A200)  and  (not A199) );
 a18300a <=( A166  and  a18299a );
 a18301a <=( a18300a  and  a18295a );
 a18304a <=( A233  and  (not A202) );
 a18308a <=( A267  and  A265 );
 a18309a <=( A234  and  a18308a );
 a18310a <=( a18309a  and  a18304a );
 a18313a <=( (not A167)  and  A170 );
 a18317a <=( (not A200)  and  (not A199) );
 a18318a <=( A166  and  a18317a );
 a18319a <=( a18318a  and  a18313a );
 a18322a <=( A233  and  (not A202) );
 a18326a <=( A267  and  A266 );
 a18327a <=( A234  and  a18326a );
 a18328a <=( a18327a  and  a18322a );
 a18331a <=( (not A167)  and  A170 );
 a18335a <=( (not A200)  and  (not A199) );
 a18336a <=( A166  and  a18335a );
 a18337a <=( a18336a  and  a18331a );
 a18340a <=( (not A232)  and  (not A202) );
 a18344a <=( A301  and  A236 );
 a18345a <=( A233  and  a18344a );
 a18346a <=( a18345a  and  a18340a );
 a18349a <=( (not A167)  and  A170 );
 a18353a <=( (not A200)  and  (not A199) );
 a18354a <=( A166  and  a18353a );
 a18355a <=( a18354a  and  a18349a );
 a18358a <=( (not A232)  and  (not A202) );
 a18362a <=( A268  and  A236 );
 a18363a <=( A233  and  a18362a );
 a18364a <=( a18363a  and  a18358a );
 a18367a <=( (not A167)  and  A170 );
 a18371a <=( (not A200)  and  (not A199) );
 a18372a <=( A166  and  a18371a );
 a18373a <=( a18372a  and  a18367a );
 a18376a <=( A232  and  (not A202) );
 a18380a <=( A301  and  A236 );
 a18381a <=( (not A233)  and  a18380a );
 a18382a <=( a18381a  and  a18376a );
 a18385a <=( (not A167)  and  A170 );
 a18389a <=( (not A200)  and  (not A199) );
 a18390a <=( A166  and  a18389a );
 a18391a <=( a18390a  and  a18385a );
 a18394a <=( A232  and  (not A202) );
 a18398a <=( A268  and  A236 );
 a18399a <=( (not A233)  and  a18398a );
 a18400a <=( a18399a  and  a18394a );
 a18403a <=( (not A201)  and  A169 );
 a18407a <=( (not A232)  and  (not A203) );
 a18408a <=( (not A202)  and  a18407a );
 a18409a <=( a18408a  and  a18403a );
 a18412a <=( A236  and  A233 );
 a18416a <=( A302  and  (not A299) );
 a18417a <=( A298  and  a18416a );
 a18418a <=( a18417a  and  a18412a );
 a18421a <=( (not A201)  and  A169 );
 a18425a <=( (not A232)  and  (not A203) );
 a18426a <=( (not A202)  and  a18425a );
 a18427a <=( a18426a  and  a18421a );
 a18430a <=( A236  and  A233 );
 a18434a <=( A302  and  A299 );
 a18435a <=( (not A298)  and  a18434a );
 a18436a <=( a18435a  and  a18430a );
 a18439a <=( (not A201)  and  A169 );
 a18443a <=( (not A232)  and  (not A203) );
 a18444a <=( (not A202)  and  a18443a );
 a18445a <=( a18444a  and  a18439a );
 a18448a <=( A236  and  A233 );
 a18452a <=( A269  and  A266 );
 a18453a <=( (not A265)  and  a18452a );
 a18454a <=( a18453a  and  a18448a );
 a18457a <=( (not A201)  and  A169 );
 a18461a <=( (not A232)  and  (not A203) );
 a18462a <=( (not A202)  and  a18461a );
 a18463a <=( a18462a  and  a18457a );
 a18466a <=( A236  and  A233 );
 a18470a <=( A269  and  (not A266) );
 a18471a <=( A265  and  a18470a );
 a18472a <=( a18471a  and  a18466a );
 a18475a <=( (not A201)  and  A169 );
 a18479a <=( A232  and  (not A203) );
 a18480a <=( (not A202)  and  a18479a );
 a18481a <=( a18480a  and  a18475a );
 a18484a <=( A236  and  (not A233) );
 a18488a <=( A302  and  (not A299) );
 a18489a <=( A298  and  a18488a );
 a18490a <=( a18489a  and  a18484a );
 a18493a <=( (not A201)  and  A169 );
 a18497a <=( A232  and  (not A203) );
 a18498a <=( (not A202)  and  a18497a );
 a18499a <=( a18498a  and  a18493a );
 a18502a <=( A236  and  (not A233) );
 a18506a <=( A302  and  A299 );
 a18507a <=( (not A298)  and  a18506a );
 a18508a <=( a18507a  and  a18502a );
 a18511a <=( (not A201)  and  A169 );
 a18515a <=( A232  and  (not A203) );
 a18516a <=( (not A202)  and  a18515a );
 a18517a <=( a18516a  and  a18511a );
 a18520a <=( A236  and  (not A233) );
 a18524a <=( A269  and  A266 );
 a18525a <=( (not A265)  and  a18524a );
 a18526a <=( a18525a  and  a18520a );
 a18529a <=( (not A201)  and  A169 );
 a18533a <=( A232  and  (not A203) );
 a18534a <=( (not A202)  and  a18533a );
 a18535a <=( a18534a  and  a18529a );
 a18538a <=( A236  and  (not A233) );
 a18542a <=( A269  and  (not A266) );
 a18543a <=( A265  and  a18542a );
 a18544a <=( a18543a  and  a18538a );
 a18547a <=( A199  and  A169 );
 a18551a <=( (not A202)  and  (not A201) );
 a18552a <=( A200  and  a18551a );
 a18553a <=( a18552a  and  a18547a );
 a18556a <=( A234  and  A232 );
 a18560a <=( A302  and  (not A299) );
 a18561a <=( A298  and  a18560a );
 a18562a <=( a18561a  and  a18556a );
 a18565a <=( A199  and  A169 );
 a18569a <=( (not A202)  and  (not A201) );
 a18570a <=( A200  and  a18569a );
 a18571a <=( a18570a  and  a18565a );
 a18574a <=( A234  and  A232 );
 a18578a <=( A302  and  A299 );
 a18579a <=( (not A298)  and  a18578a );
 a18580a <=( a18579a  and  a18574a );
 a18583a <=( A199  and  A169 );
 a18587a <=( (not A202)  and  (not A201) );
 a18588a <=( A200  and  a18587a );
 a18589a <=( a18588a  and  a18583a );
 a18592a <=( A234  and  A232 );
 a18596a <=( A269  and  A266 );
 a18597a <=( (not A265)  and  a18596a );
 a18598a <=( a18597a  and  a18592a );
 a18601a <=( A199  and  A169 );
 a18605a <=( (not A202)  and  (not A201) );
 a18606a <=( A200  and  a18605a );
 a18607a <=( a18606a  and  a18601a );
 a18610a <=( A234  and  A232 );
 a18614a <=( A269  and  (not A266) );
 a18615a <=( A265  and  a18614a );
 a18616a <=( a18615a  and  a18610a );
 a18619a <=( A199  and  A169 );
 a18623a <=( (not A202)  and  (not A201) );
 a18624a <=( A200  and  a18623a );
 a18625a <=( a18624a  and  a18619a );
 a18628a <=( A234  and  A233 );
 a18632a <=( A302  and  (not A299) );
 a18633a <=( A298  and  a18632a );
 a18634a <=( a18633a  and  a18628a );
 a18637a <=( A199  and  A169 );
 a18641a <=( (not A202)  and  (not A201) );
 a18642a <=( A200  and  a18641a );
 a18643a <=( a18642a  and  a18637a );
 a18646a <=( A234  and  A233 );
 a18650a <=( A302  and  A299 );
 a18651a <=( (not A298)  and  a18650a );
 a18652a <=( a18651a  and  a18646a );
 a18655a <=( A199  and  A169 );
 a18659a <=( (not A202)  and  (not A201) );
 a18660a <=( A200  and  a18659a );
 a18661a <=( a18660a  and  a18655a );
 a18664a <=( A234  and  A233 );
 a18668a <=( A269  and  A266 );
 a18669a <=( (not A265)  and  a18668a );
 a18670a <=( a18669a  and  a18664a );
 a18673a <=( A199  and  A169 );
 a18677a <=( (not A202)  and  (not A201) );
 a18678a <=( A200  and  a18677a );
 a18679a <=( a18678a  and  a18673a );
 a18682a <=( A234  and  A233 );
 a18686a <=( A269  and  (not A266) );
 a18687a <=( A265  and  a18686a );
 a18688a <=( a18687a  and  a18682a );
 a18691a <=( A199  and  A169 );
 a18695a <=( (not A202)  and  (not A201) );
 a18696a <=( A200  and  a18695a );
 a18697a <=( a18696a  and  a18691a );
 a18700a <=( A233  and  (not A232) );
 a18704a <=( A300  and  A299 );
 a18705a <=( A236  and  a18704a );
 a18706a <=( a18705a  and  a18700a );
 a18709a <=( A199  and  A169 );
 a18713a <=( (not A202)  and  (not A201) );
 a18714a <=( A200  and  a18713a );
 a18715a <=( a18714a  and  a18709a );
 a18718a <=( A233  and  (not A232) );
 a18722a <=( A300  and  A298 );
 a18723a <=( A236  and  a18722a );
 a18724a <=( a18723a  and  a18718a );
 a18727a <=( A199  and  A169 );
 a18731a <=( (not A202)  and  (not A201) );
 a18732a <=( A200  and  a18731a );
 a18733a <=( a18732a  and  a18727a );
 a18736a <=( A233  and  (not A232) );
 a18740a <=( A267  and  A265 );
 a18741a <=( A236  and  a18740a );
 a18742a <=( a18741a  and  a18736a );
 a18745a <=( A199  and  A169 );
 a18749a <=( (not A202)  and  (not A201) );
 a18750a <=( A200  and  a18749a );
 a18751a <=( a18750a  and  a18745a );
 a18754a <=( A233  and  (not A232) );
 a18758a <=( A267  and  A266 );
 a18759a <=( A236  and  a18758a );
 a18760a <=( a18759a  and  a18754a );
 a18763a <=( A199  and  A169 );
 a18767a <=( (not A202)  and  (not A201) );
 a18768a <=( A200  and  a18767a );
 a18769a <=( a18768a  and  a18763a );
 a18772a <=( (not A233)  and  A232 );
 a18776a <=( A300  and  A299 );
 a18777a <=( A236  and  a18776a );
 a18778a <=( a18777a  and  a18772a );
 a18781a <=( A199  and  A169 );
 a18785a <=( (not A202)  and  (not A201) );
 a18786a <=( A200  and  a18785a );
 a18787a <=( a18786a  and  a18781a );
 a18790a <=( (not A233)  and  A232 );
 a18794a <=( A300  and  A298 );
 a18795a <=( A236  and  a18794a );
 a18796a <=( a18795a  and  a18790a );
 a18799a <=( A199  and  A169 );
 a18803a <=( (not A202)  and  (not A201) );
 a18804a <=( A200  and  a18803a );
 a18805a <=( a18804a  and  a18799a );
 a18808a <=( (not A233)  and  A232 );
 a18812a <=( A267  and  A265 );
 a18813a <=( A236  and  a18812a );
 a18814a <=( a18813a  and  a18808a );
 a18817a <=( A199  and  A169 );
 a18821a <=( (not A202)  and  (not A201) );
 a18822a <=( A200  and  a18821a );
 a18823a <=( a18822a  and  a18817a );
 a18826a <=( (not A233)  and  A232 );
 a18830a <=( A267  and  A266 );
 a18831a <=( A236  and  a18830a );
 a18832a <=( a18831a  and  a18826a );
 a18835a <=( (not A199)  and  A169 );
 a18839a <=( (not A232)  and  (not A202) );
 a18840a <=( (not A200)  and  a18839a );
 a18841a <=( a18840a  and  a18835a );
 a18844a <=( A236  and  A233 );
 a18848a <=( A302  and  (not A299) );
 a18849a <=( A298  and  a18848a );
 a18850a <=( a18849a  and  a18844a );
 a18853a <=( (not A199)  and  A169 );
 a18857a <=( (not A232)  and  (not A202) );
 a18858a <=( (not A200)  and  a18857a );
 a18859a <=( a18858a  and  a18853a );
 a18862a <=( A236  and  A233 );
 a18866a <=( A302  and  A299 );
 a18867a <=( (not A298)  and  a18866a );
 a18868a <=( a18867a  and  a18862a );
 a18871a <=( (not A199)  and  A169 );
 a18875a <=( (not A232)  and  (not A202) );
 a18876a <=( (not A200)  and  a18875a );
 a18877a <=( a18876a  and  a18871a );
 a18880a <=( A236  and  A233 );
 a18884a <=( A269  and  A266 );
 a18885a <=( (not A265)  and  a18884a );
 a18886a <=( a18885a  and  a18880a );
 a18889a <=( (not A199)  and  A169 );
 a18893a <=( (not A232)  and  (not A202) );
 a18894a <=( (not A200)  and  a18893a );
 a18895a <=( a18894a  and  a18889a );
 a18898a <=( A236  and  A233 );
 a18902a <=( A269  and  (not A266) );
 a18903a <=( A265  and  a18902a );
 a18904a <=( a18903a  and  a18898a );
 a18907a <=( (not A199)  and  A169 );
 a18911a <=( A232  and  (not A202) );
 a18912a <=( (not A200)  and  a18911a );
 a18913a <=( a18912a  and  a18907a );
 a18916a <=( A236  and  (not A233) );
 a18920a <=( A302  and  (not A299) );
 a18921a <=( A298  and  a18920a );
 a18922a <=( a18921a  and  a18916a );
 a18925a <=( (not A199)  and  A169 );
 a18929a <=( A232  and  (not A202) );
 a18930a <=( (not A200)  and  a18929a );
 a18931a <=( a18930a  and  a18925a );
 a18934a <=( A236  and  (not A233) );
 a18938a <=( A302  and  A299 );
 a18939a <=( (not A298)  and  a18938a );
 a18940a <=( a18939a  and  a18934a );
 a18943a <=( (not A199)  and  A169 );
 a18947a <=( A232  and  (not A202) );
 a18948a <=( (not A200)  and  a18947a );
 a18949a <=( a18948a  and  a18943a );
 a18952a <=( A236  and  (not A233) );
 a18956a <=( A269  and  A266 );
 a18957a <=( (not A265)  and  a18956a );
 a18958a <=( a18957a  and  a18952a );
 a18961a <=( (not A199)  and  A169 );
 a18965a <=( A232  and  (not A202) );
 a18966a <=( (not A200)  and  a18965a );
 a18967a <=( a18966a  and  a18961a );
 a18970a <=( A236  and  (not A233) );
 a18974a <=( A269  and  (not A266) );
 a18975a <=( A265  and  a18974a );
 a18976a <=( a18975a  and  a18970a );
 a18979a <=( (not A167)  and  (not A169) );
 a18983a <=( (not A232)  and  A202 );
 a18984a <=( (not A166)  and  a18983a );
 a18985a <=( a18984a  and  a18979a );
 a18988a <=( A236  and  A233 );
 a18992a <=( A302  and  (not A299) );
 a18993a <=( A298  and  a18992a );
 a18994a <=( a18993a  and  a18988a );
 a18997a <=( (not A167)  and  (not A169) );
 a19001a <=( (not A232)  and  A202 );
 a19002a <=( (not A166)  and  a19001a );
 a19003a <=( a19002a  and  a18997a );
 a19006a <=( A236  and  A233 );
 a19010a <=( A302  and  A299 );
 a19011a <=( (not A298)  and  a19010a );
 a19012a <=( a19011a  and  a19006a );
 a19015a <=( (not A167)  and  (not A169) );
 a19019a <=( (not A232)  and  A202 );
 a19020a <=( (not A166)  and  a19019a );
 a19021a <=( a19020a  and  a19015a );
 a19024a <=( A236  and  A233 );
 a19028a <=( A269  and  A266 );
 a19029a <=( (not A265)  and  a19028a );
 a19030a <=( a19029a  and  a19024a );
 a19033a <=( (not A167)  and  (not A169) );
 a19037a <=( (not A232)  and  A202 );
 a19038a <=( (not A166)  and  a19037a );
 a19039a <=( a19038a  and  a19033a );
 a19042a <=( A236  and  A233 );
 a19046a <=( A269  and  (not A266) );
 a19047a <=( A265  and  a19046a );
 a19048a <=( a19047a  and  a19042a );
 a19051a <=( (not A167)  and  (not A169) );
 a19055a <=( A232  and  A202 );
 a19056a <=( (not A166)  and  a19055a );
 a19057a <=( a19056a  and  a19051a );
 a19060a <=( A236  and  (not A233) );
 a19064a <=( A302  and  (not A299) );
 a19065a <=( A298  and  a19064a );
 a19066a <=( a19065a  and  a19060a );
 a19069a <=( (not A167)  and  (not A169) );
 a19073a <=( A232  and  A202 );
 a19074a <=( (not A166)  and  a19073a );
 a19075a <=( a19074a  and  a19069a );
 a19078a <=( A236  and  (not A233) );
 a19082a <=( A302  and  A299 );
 a19083a <=( (not A298)  and  a19082a );
 a19084a <=( a19083a  and  a19078a );
 a19087a <=( (not A167)  and  (not A169) );
 a19091a <=( A232  and  A202 );
 a19092a <=( (not A166)  and  a19091a );
 a19093a <=( a19092a  and  a19087a );
 a19096a <=( A236  and  (not A233) );
 a19100a <=( A269  and  A266 );
 a19101a <=( (not A265)  and  a19100a );
 a19102a <=( a19101a  and  a19096a );
 a19105a <=( (not A167)  and  (not A169) );
 a19109a <=( A232  and  A202 );
 a19110a <=( (not A166)  and  a19109a );
 a19111a <=( a19110a  and  a19105a );
 a19114a <=( A236  and  (not A233) );
 a19118a <=( A269  and  (not A266) );
 a19119a <=( A265  and  a19118a );
 a19120a <=( a19119a  and  a19114a );
 a19123a <=( (not A167)  and  (not A169) );
 a19127a <=( A201  and  A199 );
 a19128a <=( (not A166)  and  a19127a );
 a19129a <=( a19128a  and  a19123a );
 a19132a <=( A234  and  A232 );
 a19136a <=( A302  and  (not A299) );
 a19137a <=( A298  and  a19136a );
 a19138a <=( a19137a  and  a19132a );
 a19141a <=( (not A167)  and  (not A169) );
 a19145a <=( A201  and  A199 );
 a19146a <=( (not A166)  and  a19145a );
 a19147a <=( a19146a  and  a19141a );
 a19150a <=( A234  and  A232 );
 a19154a <=( A302  and  A299 );
 a19155a <=( (not A298)  and  a19154a );
 a19156a <=( a19155a  and  a19150a );
 a19159a <=( (not A167)  and  (not A169) );
 a19163a <=( A201  and  A199 );
 a19164a <=( (not A166)  and  a19163a );
 a19165a <=( a19164a  and  a19159a );
 a19168a <=( A234  and  A232 );
 a19172a <=( A269  and  A266 );
 a19173a <=( (not A265)  and  a19172a );
 a19174a <=( a19173a  and  a19168a );
 a19177a <=( (not A167)  and  (not A169) );
 a19181a <=( A201  and  A199 );
 a19182a <=( (not A166)  and  a19181a );
 a19183a <=( a19182a  and  a19177a );
 a19186a <=( A234  and  A232 );
 a19190a <=( A269  and  (not A266) );
 a19191a <=( A265  and  a19190a );
 a19192a <=( a19191a  and  a19186a );
 a19195a <=( (not A167)  and  (not A169) );
 a19199a <=( A201  and  A199 );
 a19200a <=( (not A166)  and  a19199a );
 a19201a <=( a19200a  and  a19195a );
 a19204a <=( A234  and  A233 );
 a19208a <=( A302  and  (not A299) );
 a19209a <=( A298  and  a19208a );
 a19210a <=( a19209a  and  a19204a );
 a19213a <=( (not A167)  and  (not A169) );
 a19217a <=( A201  and  A199 );
 a19218a <=( (not A166)  and  a19217a );
 a19219a <=( a19218a  and  a19213a );
 a19222a <=( A234  and  A233 );
 a19226a <=( A302  and  A299 );
 a19227a <=( (not A298)  and  a19226a );
 a19228a <=( a19227a  and  a19222a );
 a19231a <=( (not A167)  and  (not A169) );
 a19235a <=( A201  and  A199 );
 a19236a <=( (not A166)  and  a19235a );
 a19237a <=( a19236a  and  a19231a );
 a19240a <=( A234  and  A233 );
 a19244a <=( A269  and  A266 );
 a19245a <=( (not A265)  and  a19244a );
 a19246a <=( a19245a  and  a19240a );
 a19249a <=( (not A167)  and  (not A169) );
 a19253a <=( A201  and  A199 );
 a19254a <=( (not A166)  and  a19253a );
 a19255a <=( a19254a  and  a19249a );
 a19258a <=( A234  and  A233 );
 a19262a <=( A269  and  (not A266) );
 a19263a <=( A265  and  a19262a );
 a19264a <=( a19263a  and  a19258a );
 a19267a <=( (not A167)  and  (not A169) );
 a19271a <=( A201  and  A199 );
 a19272a <=( (not A166)  and  a19271a );
 a19273a <=( a19272a  and  a19267a );
 a19276a <=( A233  and  (not A232) );
 a19280a <=( A300  and  A299 );
 a19281a <=( A236  and  a19280a );
 a19282a <=( a19281a  and  a19276a );
 a19285a <=( (not A167)  and  (not A169) );
 a19289a <=( A201  and  A199 );
 a19290a <=( (not A166)  and  a19289a );
 a19291a <=( a19290a  and  a19285a );
 a19294a <=( A233  and  (not A232) );
 a19298a <=( A300  and  A298 );
 a19299a <=( A236  and  a19298a );
 a19300a <=( a19299a  and  a19294a );
 a19303a <=( (not A167)  and  (not A169) );
 a19307a <=( A201  and  A199 );
 a19308a <=( (not A166)  and  a19307a );
 a19309a <=( a19308a  and  a19303a );
 a19312a <=( A233  and  (not A232) );
 a19316a <=( A267  and  A265 );
 a19317a <=( A236  and  a19316a );
 a19318a <=( a19317a  and  a19312a );
 a19321a <=( (not A167)  and  (not A169) );
 a19325a <=( A201  and  A199 );
 a19326a <=( (not A166)  and  a19325a );
 a19327a <=( a19326a  and  a19321a );
 a19330a <=( A233  and  (not A232) );
 a19334a <=( A267  and  A266 );
 a19335a <=( A236  and  a19334a );
 a19336a <=( a19335a  and  a19330a );
 a19339a <=( (not A167)  and  (not A169) );
 a19343a <=( A201  and  A199 );
 a19344a <=( (not A166)  and  a19343a );
 a19345a <=( a19344a  and  a19339a );
 a19348a <=( (not A233)  and  A232 );
 a19352a <=( A300  and  A299 );
 a19353a <=( A236  and  a19352a );
 a19354a <=( a19353a  and  a19348a );
 a19357a <=( (not A167)  and  (not A169) );
 a19361a <=( A201  and  A199 );
 a19362a <=( (not A166)  and  a19361a );
 a19363a <=( a19362a  and  a19357a );
 a19366a <=( (not A233)  and  A232 );
 a19370a <=( A300  and  A298 );
 a19371a <=( A236  and  a19370a );
 a19372a <=( a19371a  and  a19366a );
 a19375a <=( (not A167)  and  (not A169) );
 a19379a <=( A201  and  A199 );
 a19380a <=( (not A166)  and  a19379a );
 a19381a <=( a19380a  and  a19375a );
 a19384a <=( (not A233)  and  A232 );
 a19388a <=( A267  and  A265 );
 a19389a <=( A236  and  a19388a );
 a19390a <=( a19389a  and  a19384a );
 a19393a <=( (not A167)  and  (not A169) );
 a19397a <=( A201  and  A199 );
 a19398a <=( (not A166)  and  a19397a );
 a19399a <=( a19398a  and  a19393a );
 a19402a <=( (not A233)  and  A232 );
 a19406a <=( A267  and  A266 );
 a19407a <=( A236  and  a19406a );
 a19408a <=( a19407a  and  a19402a );
 a19411a <=( (not A167)  and  (not A169) );
 a19415a <=( A201  and  A200 );
 a19416a <=( (not A166)  and  a19415a );
 a19417a <=( a19416a  and  a19411a );
 a19420a <=( A234  and  A232 );
 a19424a <=( A302  and  (not A299) );
 a19425a <=( A298  and  a19424a );
 a19426a <=( a19425a  and  a19420a );
 a19429a <=( (not A167)  and  (not A169) );
 a19433a <=( A201  and  A200 );
 a19434a <=( (not A166)  and  a19433a );
 a19435a <=( a19434a  and  a19429a );
 a19438a <=( A234  and  A232 );
 a19442a <=( A302  and  A299 );
 a19443a <=( (not A298)  and  a19442a );
 a19444a <=( a19443a  and  a19438a );
 a19447a <=( (not A167)  and  (not A169) );
 a19451a <=( A201  and  A200 );
 a19452a <=( (not A166)  and  a19451a );
 a19453a <=( a19452a  and  a19447a );
 a19456a <=( A234  and  A232 );
 a19460a <=( A269  and  A266 );
 a19461a <=( (not A265)  and  a19460a );
 a19462a <=( a19461a  and  a19456a );
 a19465a <=( (not A167)  and  (not A169) );
 a19469a <=( A201  and  A200 );
 a19470a <=( (not A166)  and  a19469a );
 a19471a <=( a19470a  and  a19465a );
 a19474a <=( A234  and  A232 );
 a19478a <=( A269  and  (not A266) );
 a19479a <=( A265  and  a19478a );
 a19480a <=( a19479a  and  a19474a );
 a19483a <=( (not A167)  and  (not A169) );
 a19487a <=( A201  and  A200 );
 a19488a <=( (not A166)  and  a19487a );
 a19489a <=( a19488a  and  a19483a );
 a19492a <=( A234  and  A233 );
 a19496a <=( A302  and  (not A299) );
 a19497a <=( A298  and  a19496a );
 a19498a <=( a19497a  and  a19492a );
 a19501a <=( (not A167)  and  (not A169) );
 a19505a <=( A201  and  A200 );
 a19506a <=( (not A166)  and  a19505a );
 a19507a <=( a19506a  and  a19501a );
 a19510a <=( A234  and  A233 );
 a19514a <=( A302  and  A299 );
 a19515a <=( (not A298)  and  a19514a );
 a19516a <=( a19515a  and  a19510a );
 a19519a <=( (not A167)  and  (not A169) );
 a19523a <=( A201  and  A200 );
 a19524a <=( (not A166)  and  a19523a );
 a19525a <=( a19524a  and  a19519a );
 a19528a <=( A234  and  A233 );
 a19532a <=( A269  and  A266 );
 a19533a <=( (not A265)  and  a19532a );
 a19534a <=( a19533a  and  a19528a );
 a19537a <=( (not A167)  and  (not A169) );
 a19541a <=( A201  and  A200 );
 a19542a <=( (not A166)  and  a19541a );
 a19543a <=( a19542a  and  a19537a );
 a19546a <=( A234  and  A233 );
 a19550a <=( A269  and  (not A266) );
 a19551a <=( A265  and  a19550a );
 a19552a <=( a19551a  and  a19546a );
 a19555a <=( (not A167)  and  (not A169) );
 a19559a <=( A201  and  A200 );
 a19560a <=( (not A166)  and  a19559a );
 a19561a <=( a19560a  and  a19555a );
 a19564a <=( A233  and  (not A232) );
 a19568a <=( A300  and  A299 );
 a19569a <=( A236  and  a19568a );
 a19570a <=( a19569a  and  a19564a );
 a19573a <=( (not A167)  and  (not A169) );
 a19577a <=( A201  and  A200 );
 a19578a <=( (not A166)  and  a19577a );
 a19579a <=( a19578a  and  a19573a );
 a19582a <=( A233  and  (not A232) );
 a19586a <=( A300  and  A298 );
 a19587a <=( A236  and  a19586a );
 a19588a <=( a19587a  and  a19582a );
 a19591a <=( (not A167)  and  (not A169) );
 a19595a <=( A201  and  A200 );
 a19596a <=( (not A166)  and  a19595a );
 a19597a <=( a19596a  and  a19591a );
 a19600a <=( A233  and  (not A232) );
 a19604a <=( A267  and  A265 );
 a19605a <=( A236  and  a19604a );
 a19606a <=( a19605a  and  a19600a );
 a19609a <=( (not A167)  and  (not A169) );
 a19613a <=( A201  and  A200 );
 a19614a <=( (not A166)  and  a19613a );
 a19615a <=( a19614a  and  a19609a );
 a19618a <=( A233  and  (not A232) );
 a19622a <=( A267  and  A266 );
 a19623a <=( A236  and  a19622a );
 a19624a <=( a19623a  and  a19618a );
 a19627a <=( (not A167)  and  (not A169) );
 a19631a <=( A201  and  A200 );
 a19632a <=( (not A166)  and  a19631a );
 a19633a <=( a19632a  and  a19627a );
 a19636a <=( (not A233)  and  A232 );
 a19640a <=( A300  and  A299 );
 a19641a <=( A236  and  a19640a );
 a19642a <=( a19641a  and  a19636a );
 a19645a <=( (not A167)  and  (not A169) );
 a19649a <=( A201  and  A200 );
 a19650a <=( (not A166)  and  a19649a );
 a19651a <=( a19650a  and  a19645a );
 a19654a <=( (not A233)  and  A232 );
 a19658a <=( A300  and  A298 );
 a19659a <=( A236  and  a19658a );
 a19660a <=( a19659a  and  a19654a );
 a19663a <=( (not A167)  and  (not A169) );
 a19667a <=( A201  and  A200 );
 a19668a <=( (not A166)  and  a19667a );
 a19669a <=( a19668a  and  a19663a );
 a19672a <=( (not A233)  and  A232 );
 a19676a <=( A267  and  A265 );
 a19677a <=( A236  and  a19676a );
 a19678a <=( a19677a  and  a19672a );
 a19681a <=( (not A167)  and  (not A169) );
 a19685a <=( A201  and  A200 );
 a19686a <=( (not A166)  and  a19685a );
 a19687a <=( a19686a  and  a19681a );
 a19690a <=( (not A233)  and  A232 );
 a19694a <=( A267  and  A266 );
 a19695a <=( A236  and  a19694a );
 a19696a <=( a19695a  and  a19690a );
 a19699a <=( (not A167)  and  (not A169) );
 a19703a <=( A200  and  (not A199) );
 a19704a <=( (not A166)  and  a19703a );
 a19705a <=( a19704a  and  a19699a );
 a19708a <=( A235  and  A203 );
 a19712a <=( A302  and  (not A299) );
 a19713a <=( A298  and  a19712a );
 a19714a <=( a19713a  and  a19708a );
 a19717a <=( (not A167)  and  (not A169) );
 a19721a <=( A200  and  (not A199) );
 a19722a <=( (not A166)  and  a19721a );
 a19723a <=( a19722a  and  a19717a );
 a19726a <=( A235  and  A203 );
 a19730a <=( A302  and  A299 );
 a19731a <=( (not A298)  and  a19730a );
 a19732a <=( a19731a  and  a19726a );
 a19735a <=( (not A167)  and  (not A169) );
 a19739a <=( A200  and  (not A199) );
 a19740a <=( (not A166)  and  a19739a );
 a19741a <=( a19740a  and  a19735a );
 a19744a <=( A235  and  A203 );
 a19748a <=( A269  and  A266 );
 a19749a <=( (not A265)  and  a19748a );
 a19750a <=( a19749a  and  a19744a );
 a19753a <=( (not A167)  and  (not A169) );
 a19757a <=( A200  and  (not A199) );
 a19758a <=( (not A166)  and  a19757a );
 a19759a <=( a19758a  and  a19753a );
 a19762a <=( A235  and  A203 );
 a19766a <=( A269  and  (not A266) );
 a19767a <=( A265  and  a19766a );
 a19768a <=( a19767a  and  a19762a );
 a19771a <=( (not A167)  and  (not A169) );
 a19775a <=( A200  and  (not A199) );
 a19776a <=( (not A166)  and  a19775a );
 a19777a <=( a19776a  and  a19771a );
 a19780a <=( A232  and  A203 );
 a19784a <=( A300  and  A299 );
 a19785a <=( A234  and  a19784a );
 a19786a <=( a19785a  and  a19780a );
 a19789a <=( (not A167)  and  (not A169) );
 a19793a <=( A200  and  (not A199) );
 a19794a <=( (not A166)  and  a19793a );
 a19795a <=( a19794a  and  a19789a );
 a19798a <=( A232  and  A203 );
 a19802a <=( A300  and  A298 );
 a19803a <=( A234  and  a19802a );
 a19804a <=( a19803a  and  a19798a );
 a19807a <=( (not A167)  and  (not A169) );
 a19811a <=( A200  and  (not A199) );
 a19812a <=( (not A166)  and  a19811a );
 a19813a <=( a19812a  and  a19807a );
 a19816a <=( A232  and  A203 );
 a19820a <=( A267  and  A265 );
 a19821a <=( A234  and  a19820a );
 a19822a <=( a19821a  and  a19816a );
 a19825a <=( (not A167)  and  (not A169) );
 a19829a <=( A200  and  (not A199) );
 a19830a <=( (not A166)  and  a19829a );
 a19831a <=( a19830a  and  a19825a );
 a19834a <=( A232  and  A203 );
 a19838a <=( A267  and  A266 );
 a19839a <=( A234  and  a19838a );
 a19840a <=( a19839a  and  a19834a );
 a19843a <=( (not A167)  and  (not A169) );
 a19847a <=( A200  and  (not A199) );
 a19848a <=( (not A166)  and  a19847a );
 a19849a <=( a19848a  and  a19843a );
 a19852a <=( A233  and  A203 );
 a19856a <=( A300  and  A299 );
 a19857a <=( A234  and  a19856a );
 a19858a <=( a19857a  and  a19852a );
 a19861a <=( (not A167)  and  (not A169) );
 a19865a <=( A200  and  (not A199) );
 a19866a <=( (not A166)  and  a19865a );
 a19867a <=( a19866a  and  a19861a );
 a19870a <=( A233  and  A203 );
 a19874a <=( A300  and  A298 );
 a19875a <=( A234  and  a19874a );
 a19876a <=( a19875a  and  a19870a );
 a19879a <=( (not A167)  and  (not A169) );
 a19883a <=( A200  and  (not A199) );
 a19884a <=( (not A166)  and  a19883a );
 a19885a <=( a19884a  and  a19879a );
 a19888a <=( A233  and  A203 );
 a19892a <=( A267  and  A265 );
 a19893a <=( A234  and  a19892a );
 a19894a <=( a19893a  and  a19888a );
 a19897a <=( (not A167)  and  (not A169) );
 a19901a <=( A200  and  (not A199) );
 a19902a <=( (not A166)  and  a19901a );
 a19903a <=( a19902a  and  a19897a );
 a19906a <=( A233  and  A203 );
 a19910a <=( A267  and  A266 );
 a19911a <=( A234  and  a19910a );
 a19912a <=( a19911a  and  a19906a );
 a19915a <=( (not A167)  and  (not A169) );
 a19919a <=( A200  and  (not A199) );
 a19920a <=( (not A166)  and  a19919a );
 a19921a <=( a19920a  and  a19915a );
 a19924a <=( (not A232)  and  A203 );
 a19928a <=( A301  and  A236 );
 a19929a <=( A233  and  a19928a );
 a19930a <=( a19929a  and  a19924a );
 a19933a <=( (not A167)  and  (not A169) );
 a19937a <=( A200  and  (not A199) );
 a19938a <=( (not A166)  and  a19937a );
 a19939a <=( a19938a  and  a19933a );
 a19942a <=( (not A232)  and  A203 );
 a19946a <=( A268  and  A236 );
 a19947a <=( A233  and  a19946a );
 a19948a <=( a19947a  and  a19942a );
 a19951a <=( (not A167)  and  (not A169) );
 a19955a <=( A200  and  (not A199) );
 a19956a <=( (not A166)  and  a19955a );
 a19957a <=( a19956a  and  a19951a );
 a19960a <=( A232  and  A203 );
 a19964a <=( A301  and  A236 );
 a19965a <=( (not A233)  and  a19964a );
 a19966a <=( a19965a  and  a19960a );
 a19969a <=( (not A167)  and  (not A169) );
 a19973a <=( A200  and  (not A199) );
 a19974a <=( (not A166)  and  a19973a );
 a19975a <=( a19974a  and  a19969a );
 a19978a <=( A232  and  A203 );
 a19982a <=( A268  and  A236 );
 a19983a <=( (not A233)  and  a19982a );
 a19984a <=( a19983a  and  a19978a );
 a19987a <=( (not A167)  and  (not A169) );
 a19991a <=( (not A200)  and  A199 );
 a19992a <=( (not A166)  and  a19991a );
 a19993a <=( a19992a  and  a19987a );
 a19996a <=( A235  and  A203 );
 a20000a <=( A302  and  (not A299) );
 a20001a <=( A298  and  a20000a );
 a20002a <=( a20001a  and  a19996a );
 a20005a <=( (not A167)  and  (not A169) );
 a20009a <=( (not A200)  and  A199 );
 a20010a <=( (not A166)  and  a20009a );
 a20011a <=( a20010a  and  a20005a );
 a20014a <=( A235  and  A203 );
 a20018a <=( A302  and  A299 );
 a20019a <=( (not A298)  and  a20018a );
 a20020a <=( a20019a  and  a20014a );
 a20023a <=( (not A167)  and  (not A169) );
 a20027a <=( (not A200)  and  A199 );
 a20028a <=( (not A166)  and  a20027a );
 a20029a <=( a20028a  and  a20023a );
 a20032a <=( A235  and  A203 );
 a20036a <=( A269  and  A266 );
 a20037a <=( (not A265)  and  a20036a );
 a20038a <=( a20037a  and  a20032a );
 a20041a <=( (not A167)  and  (not A169) );
 a20045a <=( (not A200)  and  A199 );
 a20046a <=( (not A166)  and  a20045a );
 a20047a <=( a20046a  and  a20041a );
 a20050a <=( A235  and  A203 );
 a20054a <=( A269  and  (not A266) );
 a20055a <=( A265  and  a20054a );
 a20056a <=( a20055a  and  a20050a );
 a20059a <=( (not A167)  and  (not A169) );
 a20063a <=( (not A200)  and  A199 );
 a20064a <=( (not A166)  and  a20063a );
 a20065a <=( a20064a  and  a20059a );
 a20068a <=( A232  and  A203 );
 a20072a <=( A300  and  A299 );
 a20073a <=( A234  and  a20072a );
 a20074a <=( a20073a  and  a20068a );
 a20077a <=( (not A167)  and  (not A169) );
 a20081a <=( (not A200)  and  A199 );
 a20082a <=( (not A166)  and  a20081a );
 a20083a <=( a20082a  and  a20077a );
 a20086a <=( A232  and  A203 );
 a20090a <=( A300  and  A298 );
 a20091a <=( A234  and  a20090a );
 a20092a <=( a20091a  and  a20086a );
 a20095a <=( (not A167)  and  (not A169) );
 a20099a <=( (not A200)  and  A199 );
 a20100a <=( (not A166)  and  a20099a );
 a20101a <=( a20100a  and  a20095a );
 a20104a <=( A232  and  A203 );
 a20108a <=( A267  and  A265 );
 a20109a <=( A234  and  a20108a );
 a20110a <=( a20109a  and  a20104a );
 a20113a <=( (not A167)  and  (not A169) );
 a20117a <=( (not A200)  and  A199 );
 a20118a <=( (not A166)  and  a20117a );
 a20119a <=( a20118a  and  a20113a );
 a20122a <=( A232  and  A203 );
 a20126a <=( A267  and  A266 );
 a20127a <=( A234  and  a20126a );
 a20128a <=( a20127a  and  a20122a );
 a20131a <=( (not A167)  and  (not A169) );
 a20135a <=( (not A200)  and  A199 );
 a20136a <=( (not A166)  and  a20135a );
 a20137a <=( a20136a  and  a20131a );
 a20140a <=( A233  and  A203 );
 a20144a <=( A300  and  A299 );
 a20145a <=( A234  and  a20144a );
 a20146a <=( a20145a  and  a20140a );
 a20149a <=( (not A167)  and  (not A169) );
 a20153a <=( (not A200)  and  A199 );
 a20154a <=( (not A166)  and  a20153a );
 a20155a <=( a20154a  and  a20149a );
 a20158a <=( A233  and  A203 );
 a20162a <=( A300  and  A298 );
 a20163a <=( A234  and  a20162a );
 a20164a <=( a20163a  and  a20158a );
 a20167a <=( (not A167)  and  (not A169) );
 a20171a <=( (not A200)  and  A199 );
 a20172a <=( (not A166)  and  a20171a );
 a20173a <=( a20172a  and  a20167a );
 a20176a <=( A233  and  A203 );
 a20180a <=( A267  and  A265 );
 a20181a <=( A234  and  a20180a );
 a20182a <=( a20181a  and  a20176a );
 a20185a <=( (not A167)  and  (not A169) );
 a20189a <=( (not A200)  and  A199 );
 a20190a <=( (not A166)  and  a20189a );
 a20191a <=( a20190a  and  a20185a );
 a20194a <=( A233  and  A203 );
 a20198a <=( A267  and  A266 );
 a20199a <=( A234  and  a20198a );
 a20200a <=( a20199a  and  a20194a );
 a20203a <=( (not A167)  and  (not A169) );
 a20207a <=( (not A200)  and  A199 );
 a20208a <=( (not A166)  and  a20207a );
 a20209a <=( a20208a  and  a20203a );
 a20212a <=( (not A232)  and  A203 );
 a20216a <=( A301  and  A236 );
 a20217a <=( A233  and  a20216a );
 a20218a <=( a20217a  and  a20212a );
 a20221a <=( (not A167)  and  (not A169) );
 a20225a <=( (not A200)  and  A199 );
 a20226a <=( (not A166)  and  a20225a );
 a20227a <=( a20226a  and  a20221a );
 a20230a <=( (not A232)  and  A203 );
 a20234a <=( A268  and  A236 );
 a20235a <=( A233  and  a20234a );
 a20236a <=( a20235a  and  a20230a );
 a20239a <=( (not A167)  and  (not A169) );
 a20243a <=( (not A200)  and  A199 );
 a20244a <=( (not A166)  and  a20243a );
 a20245a <=( a20244a  and  a20239a );
 a20248a <=( A232  and  A203 );
 a20252a <=( A301  and  A236 );
 a20253a <=( (not A233)  and  a20252a );
 a20254a <=( a20253a  and  a20248a );
 a20257a <=( (not A167)  and  (not A169) );
 a20261a <=( (not A200)  and  A199 );
 a20262a <=( (not A166)  and  a20261a );
 a20263a <=( a20262a  and  a20257a );
 a20266a <=( A232  and  A203 );
 a20270a <=( A268  and  A236 );
 a20271a <=( (not A233)  and  a20270a );
 a20272a <=( a20271a  and  a20266a );
 a20275a <=( (not A168)  and  (not A169) );
 a20279a <=( A202  and  A166 );
 a20280a <=( A167  and  a20279a );
 a20281a <=( a20280a  and  a20275a );
 a20284a <=( A234  and  A232 );
 a20288a <=( A302  and  (not A299) );
 a20289a <=( A298  and  a20288a );
 a20290a <=( a20289a  and  a20284a );
 a20293a <=( (not A168)  and  (not A169) );
 a20297a <=( A202  and  A166 );
 a20298a <=( A167  and  a20297a );
 a20299a <=( a20298a  and  a20293a );
 a20302a <=( A234  and  A232 );
 a20306a <=( A302  and  A299 );
 a20307a <=( (not A298)  and  a20306a );
 a20308a <=( a20307a  and  a20302a );
 a20311a <=( (not A168)  and  (not A169) );
 a20315a <=( A202  and  A166 );
 a20316a <=( A167  and  a20315a );
 a20317a <=( a20316a  and  a20311a );
 a20320a <=( A234  and  A232 );
 a20324a <=( A269  and  A266 );
 a20325a <=( (not A265)  and  a20324a );
 a20326a <=( a20325a  and  a20320a );
 a20329a <=( (not A168)  and  (not A169) );
 a20333a <=( A202  and  A166 );
 a20334a <=( A167  and  a20333a );
 a20335a <=( a20334a  and  a20329a );
 a20338a <=( A234  and  A232 );
 a20342a <=( A269  and  (not A266) );
 a20343a <=( A265  and  a20342a );
 a20344a <=( a20343a  and  a20338a );
 a20347a <=( (not A168)  and  (not A169) );
 a20351a <=( A202  and  A166 );
 a20352a <=( A167  and  a20351a );
 a20353a <=( a20352a  and  a20347a );
 a20356a <=( A234  and  A233 );
 a20360a <=( A302  and  (not A299) );
 a20361a <=( A298  and  a20360a );
 a20362a <=( a20361a  and  a20356a );
 a20365a <=( (not A168)  and  (not A169) );
 a20369a <=( A202  and  A166 );
 a20370a <=( A167  and  a20369a );
 a20371a <=( a20370a  and  a20365a );
 a20374a <=( A234  and  A233 );
 a20378a <=( A302  and  A299 );
 a20379a <=( (not A298)  and  a20378a );
 a20380a <=( a20379a  and  a20374a );
 a20383a <=( (not A168)  and  (not A169) );
 a20387a <=( A202  and  A166 );
 a20388a <=( A167  and  a20387a );
 a20389a <=( a20388a  and  a20383a );
 a20392a <=( A234  and  A233 );
 a20396a <=( A269  and  A266 );
 a20397a <=( (not A265)  and  a20396a );
 a20398a <=( a20397a  and  a20392a );
 a20401a <=( (not A168)  and  (not A169) );
 a20405a <=( A202  and  A166 );
 a20406a <=( A167  and  a20405a );
 a20407a <=( a20406a  and  a20401a );
 a20410a <=( A234  and  A233 );
 a20414a <=( A269  and  (not A266) );
 a20415a <=( A265  and  a20414a );
 a20416a <=( a20415a  and  a20410a );
 a20419a <=( (not A168)  and  (not A169) );
 a20423a <=( A202  and  A166 );
 a20424a <=( A167  and  a20423a );
 a20425a <=( a20424a  and  a20419a );
 a20428a <=( A233  and  (not A232) );
 a20432a <=( A300  and  A299 );
 a20433a <=( A236  and  a20432a );
 a20434a <=( a20433a  and  a20428a );
 a20437a <=( (not A168)  and  (not A169) );
 a20441a <=( A202  and  A166 );
 a20442a <=( A167  and  a20441a );
 a20443a <=( a20442a  and  a20437a );
 a20446a <=( A233  and  (not A232) );
 a20450a <=( A300  and  A298 );
 a20451a <=( A236  and  a20450a );
 a20452a <=( a20451a  and  a20446a );
 a20455a <=( (not A168)  and  (not A169) );
 a20459a <=( A202  and  A166 );
 a20460a <=( A167  and  a20459a );
 a20461a <=( a20460a  and  a20455a );
 a20464a <=( A233  and  (not A232) );
 a20468a <=( A267  and  A265 );
 a20469a <=( A236  and  a20468a );
 a20470a <=( a20469a  and  a20464a );
 a20473a <=( (not A168)  and  (not A169) );
 a20477a <=( A202  and  A166 );
 a20478a <=( A167  and  a20477a );
 a20479a <=( a20478a  and  a20473a );
 a20482a <=( A233  and  (not A232) );
 a20486a <=( A267  and  A266 );
 a20487a <=( A236  and  a20486a );
 a20488a <=( a20487a  and  a20482a );
 a20491a <=( (not A168)  and  (not A169) );
 a20495a <=( A202  and  A166 );
 a20496a <=( A167  and  a20495a );
 a20497a <=( a20496a  and  a20491a );
 a20500a <=( (not A233)  and  A232 );
 a20504a <=( A300  and  A299 );
 a20505a <=( A236  and  a20504a );
 a20506a <=( a20505a  and  a20500a );
 a20509a <=( (not A168)  and  (not A169) );
 a20513a <=( A202  and  A166 );
 a20514a <=( A167  and  a20513a );
 a20515a <=( a20514a  and  a20509a );
 a20518a <=( (not A233)  and  A232 );
 a20522a <=( A300  and  A298 );
 a20523a <=( A236  and  a20522a );
 a20524a <=( a20523a  and  a20518a );
 a20527a <=( (not A168)  and  (not A169) );
 a20531a <=( A202  and  A166 );
 a20532a <=( A167  and  a20531a );
 a20533a <=( a20532a  and  a20527a );
 a20536a <=( (not A233)  and  A232 );
 a20540a <=( A267  and  A265 );
 a20541a <=( A236  and  a20540a );
 a20542a <=( a20541a  and  a20536a );
 a20545a <=( (not A168)  and  (not A169) );
 a20549a <=( A202  and  A166 );
 a20550a <=( A167  and  a20549a );
 a20551a <=( a20550a  and  a20545a );
 a20554a <=( (not A233)  and  A232 );
 a20558a <=( A267  and  A266 );
 a20559a <=( A236  and  a20558a );
 a20560a <=( a20559a  and  a20554a );
 a20563a <=( (not A168)  and  (not A169) );
 a20567a <=( A199  and  A166 );
 a20568a <=( A167  and  a20567a );
 a20569a <=( a20568a  and  a20563a );
 a20572a <=( A235  and  A201 );
 a20576a <=( A302  and  (not A299) );
 a20577a <=( A298  and  a20576a );
 a20578a <=( a20577a  and  a20572a );
 a20581a <=( (not A168)  and  (not A169) );
 a20585a <=( A199  and  A166 );
 a20586a <=( A167  and  a20585a );
 a20587a <=( a20586a  and  a20581a );
 a20590a <=( A235  and  A201 );
 a20594a <=( A302  and  A299 );
 a20595a <=( (not A298)  and  a20594a );
 a20596a <=( a20595a  and  a20590a );
 a20599a <=( (not A168)  and  (not A169) );
 a20603a <=( A199  and  A166 );
 a20604a <=( A167  and  a20603a );
 a20605a <=( a20604a  and  a20599a );
 a20608a <=( A235  and  A201 );
 a20612a <=( A269  and  A266 );
 a20613a <=( (not A265)  and  a20612a );
 a20614a <=( a20613a  and  a20608a );
 a20617a <=( (not A168)  and  (not A169) );
 a20621a <=( A199  and  A166 );
 a20622a <=( A167  and  a20621a );
 a20623a <=( a20622a  and  a20617a );
 a20626a <=( A235  and  A201 );
 a20630a <=( A269  and  (not A266) );
 a20631a <=( A265  and  a20630a );
 a20632a <=( a20631a  and  a20626a );
 a20635a <=( (not A168)  and  (not A169) );
 a20639a <=( A199  and  A166 );
 a20640a <=( A167  and  a20639a );
 a20641a <=( a20640a  and  a20635a );
 a20644a <=( A232  and  A201 );
 a20648a <=( A300  and  A299 );
 a20649a <=( A234  and  a20648a );
 a20650a <=( a20649a  and  a20644a );
 a20653a <=( (not A168)  and  (not A169) );
 a20657a <=( A199  and  A166 );
 a20658a <=( A167  and  a20657a );
 a20659a <=( a20658a  and  a20653a );
 a20662a <=( A232  and  A201 );
 a20666a <=( A300  and  A298 );
 a20667a <=( A234  and  a20666a );
 a20668a <=( a20667a  and  a20662a );
 a20671a <=( (not A168)  and  (not A169) );
 a20675a <=( A199  and  A166 );
 a20676a <=( A167  and  a20675a );
 a20677a <=( a20676a  and  a20671a );
 a20680a <=( A232  and  A201 );
 a20684a <=( A267  and  A265 );
 a20685a <=( A234  and  a20684a );
 a20686a <=( a20685a  and  a20680a );
 a20689a <=( (not A168)  and  (not A169) );
 a20693a <=( A199  and  A166 );
 a20694a <=( A167  and  a20693a );
 a20695a <=( a20694a  and  a20689a );
 a20698a <=( A232  and  A201 );
 a20702a <=( A267  and  A266 );
 a20703a <=( A234  and  a20702a );
 a20704a <=( a20703a  and  a20698a );
 a20707a <=( (not A168)  and  (not A169) );
 a20711a <=( A199  and  A166 );
 a20712a <=( A167  and  a20711a );
 a20713a <=( a20712a  and  a20707a );
 a20716a <=( A233  and  A201 );
 a20720a <=( A300  and  A299 );
 a20721a <=( A234  and  a20720a );
 a20722a <=( a20721a  and  a20716a );
 a20725a <=( (not A168)  and  (not A169) );
 a20729a <=( A199  and  A166 );
 a20730a <=( A167  and  a20729a );
 a20731a <=( a20730a  and  a20725a );
 a20734a <=( A233  and  A201 );
 a20738a <=( A300  and  A298 );
 a20739a <=( A234  and  a20738a );
 a20740a <=( a20739a  and  a20734a );
 a20743a <=( (not A168)  and  (not A169) );
 a20747a <=( A199  and  A166 );
 a20748a <=( A167  and  a20747a );
 a20749a <=( a20748a  and  a20743a );
 a20752a <=( A233  and  A201 );
 a20756a <=( A267  and  A265 );
 a20757a <=( A234  and  a20756a );
 a20758a <=( a20757a  and  a20752a );
 a20761a <=( (not A168)  and  (not A169) );
 a20765a <=( A199  and  A166 );
 a20766a <=( A167  and  a20765a );
 a20767a <=( a20766a  and  a20761a );
 a20770a <=( A233  and  A201 );
 a20774a <=( A267  and  A266 );
 a20775a <=( A234  and  a20774a );
 a20776a <=( a20775a  and  a20770a );
 a20779a <=( (not A168)  and  (not A169) );
 a20783a <=( A199  and  A166 );
 a20784a <=( A167  and  a20783a );
 a20785a <=( a20784a  and  a20779a );
 a20788a <=( (not A232)  and  A201 );
 a20792a <=( A301  and  A236 );
 a20793a <=( A233  and  a20792a );
 a20794a <=( a20793a  and  a20788a );
 a20797a <=( (not A168)  and  (not A169) );
 a20801a <=( A199  and  A166 );
 a20802a <=( A167  and  a20801a );
 a20803a <=( a20802a  and  a20797a );
 a20806a <=( (not A232)  and  A201 );
 a20810a <=( A268  and  A236 );
 a20811a <=( A233  and  a20810a );
 a20812a <=( a20811a  and  a20806a );
 a20815a <=( (not A168)  and  (not A169) );
 a20819a <=( A199  and  A166 );
 a20820a <=( A167  and  a20819a );
 a20821a <=( a20820a  and  a20815a );
 a20824a <=( A232  and  A201 );
 a20828a <=( A301  and  A236 );
 a20829a <=( (not A233)  and  a20828a );
 a20830a <=( a20829a  and  a20824a );
 a20833a <=( (not A168)  and  (not A169) );
 a20837a <=( A199  and  A166 );
 a20838a <=( A167  and  a20837a );
 a20839a <=( a20838a  and  a20833a );
 a20842a <=( A232  and  A201 );
 a20846a <=( A268  and  A236 );
 a20847a <=( (not A233)  and  a20846a );
 a20848a <=( a20847a  and  a20842a );
 a20851a <=( (not A168)  and  (not A169) );
 a20855a <=( A200  and  A166 );
 a20856a <=( A167  and  a20855a );
 a20857a <=( a20856a  and  a20851a );
 a20860a <=( A235  and  A201 );
 a20864a <=( A302  and  (not A299) );
 a20865a <=( A298  and  a20864a );
 a20866a <=( a20865a  and  a20860a );
 a20869a <=( (not A168)  and  (not A169) );
 a20873a <=( A200  and  A166 );
 a20874a <=( A167  and  a20873a );
 a20875a <=( a20874a  and  a20869a );
 a20878a <=( A235  and  A201 );
 a20882a <=( A302  and  A299 );
 a20883a <=( (not A298)  and  a20882a );
 a20884a <=( a20883a  and  a20878a );
 a20887a <=( (not A168)  and  (not A169) );
 a20891a <=( A200  and  A166 );
 a20892a <=( A167  and  a20891a );
 a20893a <=( a20892a  and  a20887a );
 a20896a <=( A235  and  A201 );
 a20900a <=( A269  and  A266 );
 a20901a <=( (not A265)  and  a20900a );
 a20902a <=( a20901a  and  a20896a );
 a20905a <=( (not A168)  and  (not A169) );
 a20909a <=( A200  and  A166 );
 a20910a <=( A167  and  a20909a );
 a20911a <=( a20910a  and  a20905a );
 a20914a <=( A235  and  A201 );
 a20918a <=( A269  and  (not A266) );
 a20919a <=( A265  and  a20918a );
 a20920a <=( a20919a  and  a20914a );
 a20923a <=( (not A168)  and  (not A169) );
 a20927a <=( A200  and  A166 );
 a20928a <=( A167  and  a20927a );
 a20929a <=( a20928a  and  a20923a );
 a20932a <=( A232  and  A201 );
 a20936a <=( A300  and  A299 );
 a20937a <=( A234  and  a20936a );
 a20938a <=( a20937a  and  a20932a );
 a20941a <=( (not A168)  and  (not A169) );
 a20945a <=( A200  and  A166 );
 a20946a <=( A167  and  a20945a );
 a20947a <=( a20946a  and  a20941a );
 a20950a <=( A232  and  A201 );
 a20954a <=( A300  and  A298 );
 a20955a <=( A234  and  a20954a );
 a20956a <=( a20955a  and  a20950a );
 a20959a <=( (not A168)  and  (not A169) );
 a20963a <=( A200  and  A166 );
 a20964a <=( A167  and  a20963a );
 a20965a <=( a20964a  and  a20959a );
 a20968a <=( A232  and  A201 );
 a20972a <=( A267  and  A265 );
 a20973a <=( A234  and  a20972a );
 a20974a <=( a20973a  and  a20968a );
 a20977a <=( (not A168)  and  (not A169) );
 a20981a <=( A200  and  A166 );
 a20982a <=( A167  and  a20981a );
 a20983a <=( a20982a  and  a20977a );
 a20986a <=( A232  and  A201 );
 a20990a <=( A267  and  A266 );
 a20991a <=( A234  and  a20990a );
 a20992a <=( a20991a  and  a20986a );
 a20995a <=( (not A168)  and  (not A169) );
 a20999a <=( A200  and  A166 );
 a21000a <=( A167  and  a20999a );
 a21001a <=( a21000a  and  a20995a );
 a21004a <=( A233  and  A201 );
 a21008a <=( A300  and  A299 );
 a21009a <=( A234  and  a21008a );
 a21010a <=( a21009a  and  a21004a );
 a21013a <=( (not A168)  and  (not A169) );
 a21017a <=( A200  and  A166 );
 a21018a <=( A167  and  a21017a );
 a21019a <=( a21018a  and  a21013a );
 a21022a <=( A233  and  A201 );
 a21026a <=( A300  and  A298 );
 a21027a <=( A234  and  a21026a );
 a21028a <=( a21027a  and  a21022a );
 a21031a <=( (not A168)  and  (not A169) );
 a21035a <=( A200  and  A166 );
 a21036a <=( A167  and  a21035a );
 a21037a <=( a21036a  and  a21031a );
 a21040a <=( A233  and  A201 );
 a21044a <=( A267  and  A265 );
 a21045a <=( A234  and  a21044a );
 a21046a <=( a21045a  and  a21040a );
 a21049a <=( (not A168)  and  (not A169) );
 a21053a <=( A200  and  A166 );
 a21054a <=( A167  and  a21053a );
 a21055a <=( a21054a  and  a21049a );
 a21058a <=( A233  and  A201 );
 a21062a <=( A267  and  A266 );
 a21063a <=( A234  and  a21062a );
 a21064a <=( a21063a  and  a21058a );
 a21067a <=( (not A168)  and  (not A169) );
 a21071a <=( A200  and  A166 );
 a21072a <=( A167  and  a21071a );
 a21073a <=( a21072a  and  a21067a );
 a21076a <=( (not A232)  and  A201 );
 a21080a <=( A301  and  A236 );
 a21081a <=( A233  and  a21080a );
 a21082a <=( a21081a  and  a21076a );
 a21085a <=( (not A168)  and  (not A169) );
 a21089a <=( A200  and  A166 );
 a21090a <=( A167  and  a21089a );
 a21091a <=( a21090a  and  a21085a );
 a21094a <=( (not A232)  and  A201 );
 a21098a <=( A268  and  A236 );
 a21099a <=( A233  and  a21098a );
 a21100a <=( a21099a  and  a21094a );
 a21103a <=( (not A168)  and  (not A169) );
 a21107a <=( A200  and  A166 );
 a21108a <=( A167  and  a21107a );
 a21109a <=( a21108a  and  a21103a );
 a21112a <=( A232  and  A201 );
 a21116a <=( A301  and  A236 );
 a21117a <=( (not A233)  and  a21116a );
 a21118a <=( a21117a  and  a21112a );
 a21121a <=( (not A168)  and  (not A169) );
 a21125a <=( A200  and  A166 );
 a21126a <=( A167  and  a21125a );
 a21127a <=( a21126a  and  a21121a );
 a21130a <=( A232  and  A201 );
 a21134a <=( A268  and  A236 );
 a21135a <=( (not A233)  and  a21134a );
 a21136a <=( a21135a  and  a21130a );
 a21139a <=( (not A168)  and  (not A169) );
 a21143a <=( (not A199)  and  A166 );
 a21144a <=( A167  and  a21143a );
 a21145a <=( a21144a  and  a21139a );
 a21148a <=( A203  and  A200 );
 a21152a <=( A300  and  A299 );
 a21153a <=( A235  and  a21152a );
 a21154a <=( a21153a  and  a21148a );
 a21157a <=( (not A168)  and  (not A169) );
 a21161a <=( (not A199)  and  A166 );
 a21162a <=( A167  and  a21161a );
 a21163a <=( a21162a  and  a21157a );
 a21166a <=( A203  and  A200 );
 a21170a <=( A300  and  A298 );
 a21171a <=( A235  and  a21170a );
 a21172a <=( a21171a  and  a21166a );
 a21175a <=( (not A168)  and  (not A169) );
 a21179a <=( (not A199)  and  A166 );
 a21180a <=( A167  and  a21179a );
 a21181a <=( a21180a  and  a21175a );
 a21184a <=( A203  and  A200 );
 a21188a <=( A267  and  A265 );
 a21189a <=( A235  and  a21188a );
 a21190a <=( a21189a  and  a21184a );
 a21193a <=( (not A168)  and  (not A169) );
 a21197a <=( (not A199)  and  A166 );
 a21198a <=( A167  and  a21197a );
 a21199a <=( a21198a  and  a21193a );
 a21202a <=( A203  and  A200 );
 a21206a <=( A267  and  A266 );
 a21207a <=( A235  and  a21206a );
 a21208a <=( a21207a  and  a21202a );
 a21211a <=( (not A168)  and  (not A169) );
 a21215a <=( (not A199)  and  A166 );
 a21216a <=( A167  and  a21215a );
 a21217a <=( a21216a  and  a21211a );
 a21220a <=( A203  and  A200 );
 a21224a <=( A301  and  A234 );
 a21225a <=( A232  and  a21224a );
 a21226a <=( a21225a  and  a21220a );
 a21229a <=( (not A168)  and  (not A169) );
 a21233a <=( (not A199)  and  A166 );
 a21234a <=( A167  and  a21233a );
 a21235a <=( a21234a  and  a21229a );
 a21238a <=( A203  and  A200 );
 a21242a <=( A268  and  A234 );
 a21243a <=( A232  and  a21242a );
 a21244a <=( a21243a  and  a21238a );
 a21247a <=( (not A168)  and  (not A169) );
 a21251a <=( (not A199)  and  A166 );
 a21252a <=( A167  and  a21251a );
 a21253a <=( a21252a  and  a21247a );
 a21256a <=( A203  and  A200 );
 a21260a <=( A301  and  A234 );
 a21261a <=( A233  and  a21260a );
 a21262a <=( a21261a  and  a21256a );
 a21265a <=( (not A168)  and  (not A169) );
 a21269a <=( (not A199)  and  A166 );
 a21270a <=( A167  and  a21269a );
 a21271a <=( a21270a  and  a21265a );
 a21274a <=( A203  and  A200 );
 a21278a <=( A268  and  A234 );
 a21279a <=( A233  and  a21278a );
 a21280a <=( a21279a  and  a21274a );
 a21283a <=( (not A168)  and  (not A169) );
 a21287a <=( A199  and  A166 );
 a21288a <=( A167  and  a21287a );
 a21289a <=( a21288a  and  a21283a );
 a21292a <=( A203  and  (not A200) );
 a21296a <=( A300  and  A299 );
 a21297a <=( A235  and  a21296a );
 a21298a <=( a21297a  and  a21292a );
 a21301a <=( (not A168)  and  (not A169) );
 a21305a <=( A199  and  A166 );
 a21306a <=( A167  and  a21305a );
 a21307a <=( a21306a  and  a21301a );
 a21310a <=( A203  and  (not A200) );
 a21314a <=( A300  and  A298 );
 a21315a <=( A235  and  a21314a );
 a21316a <=( a21315a  and  a21310a );
 a21319a <=( (not A168)  and  (not A169) );
 a21323a <=( A199  and  A166 );
 a21324a <=( A167  and  a21323a );
 a21325a <=( a21324a  and  a21319a );
 a21328a <=( A203  and  (not A200) );
 a21332a <=( A267  and  A265 );
 a21333a <=( A235  and  a21332a );
 a21334a <=( a21333a  and  a21328a );
 a21337a <=( (not A168)  and  (not A169) );
 a21341a <=( A199  and  A166 );
 a21342a <=( A167  and  a21341a );
 a21343a <=( a21342a  and  a21337a );
 a21346a <=( A203  and  (not A200) );
 a21350a <=( A267  and  A266 );
 a21351a <=( A235  and  a21350a );
 a21352a <=( a21351a  and  a21346a );
 a21355a <=( (not A168)  and  (not A169) );
 a21359a <=( A199  and  A166 );
 a21360a <=( A167  and  a21359a );
 a21361a <=( a21360a  and  a21355a );
 a21364a <=( A203  and  (not A200) );
 a21368a <=( A301  and  A234 );
 a21369a <=( A232  and  a21368a );
 a21370a <=( a21369a  and  a21364a );
 a21373a <=( (not A168)  and  (not A169) );
 a21377a <=( A199  and  A166 );
 a21378a <=( A167  and  a21377a );
 a21379a <=( a21378a  and  a21373a );
 a21382a <=( A203  and  (not A200) );
 a21386a <=( A268  and  A234 );
 a21387a <=( A232  and  a21386a );
 a21388a <=( a21387a  and  a21382a );
 a21391a <=( (not A168)  and  (not A169) );
 a21395a <=( A199  and  A166 );
 a21396a <=( A167  and  a21395a );
 a21397a <=( a21396a  and  a21391a );
 a21400a <=( A203  and  (not A200) );
 a21404a <=( A301  and  A234 );
 a21405a <=( A233  and  a21404a );
 a21406a <=( a21405a  and  a21400a );
 a21409a <=( (not A168)  and  (not A169) );
 a21413a <=( A199  and  A166 );
 a21414a <=( A167  and  a21413a );
 a21415a <=( a21414a  and  a21409a );
 a21418a <=( A203  and  (not A200) );
 a21422a <=( A268  and  A234 );
 a21423a <=( A233  and  a21422a );
 a21424a <=( a21423a  and  a21418a );
 a21427a <=( (not A169)  and  (not A170) );
 a21431a <=( (not A232)  and  A202 );
 a21432a <=( (not A168)  and  a21431a );
 a21433a <=( a21432a  and  a21427a );
 a21436a <=( A236  and  A233 );
 a21440a <=( A302  and  (not A299) );
 a21441a <=( A298  and  a21440a );
 a21442a <=( a21441a  and  a21436a );
 a21445a <=( (not A169)  and  (not A170) );
 a21449a <=( (not A232)  and  A202 );
 a21450a <=( (not A168)  and  a21449a );
 a21451a <=( a21450a  and  a21445a );
 a21454a <=( A236  and  A233 );
 a21458a <=( A302  and  A299 );
 a21459a <=( (not A298)  and  a21458a );
 a21460a <=( a21459a  and  a21454a );
 a21463a <=( (not A169)  and  (not A170) );
 a21467a <=( (not A232)  and  A202 );
 a21468a <=( (not A168)  and  a21467a );
 a21469a <=( a21468a  and  a21463a );
 a21472a <=( A236  and  A233 );
 a21476a <=( A269  and  A266 );
 a21477a <=( (not A265)  and  a21476a );
 a21478a <=( a21477a  and  a21472a );
 a21481a <=( (not A169)  and  (not A170) );
 a21485a <=( (not A232)  and  A202 );
 a21486a <=( (not A168)  and  a21485a );
 a21487a <=( a21486a  and  a21481a );
 a21490a <=( A236  and  A233 );
 a21494a <=( A269  and  (not A266) );
 a21495a <=( A265  and  a21494a );
 a21496a <=( a21495a  and  a21490a );
 a21499a <=( (not A169)  and  (not A170) );
 a21503a <=( A232  and  A202 );
 a21504a <=( (not A168)  and  a21503a );
 a21505a <=( a21504a  and  a21499a );
 a21508a <=( A236  and  (not A233) );
 a21512a <=( A302  and  (not A299) );
 a21513a <=( A298  and  a21512a );
 a21514a <=( a21513a  and  a21508a );
 a21517a <=( (not A169)  and  (not A170) );
 a21521a <=( A232  and  A202 );
 a21522a <=( (not A168)  and  a21521a );
 a21523a <=( a21522a  and  a21517a );
 a21526a <=( A236  and  (not A233) );
 a21530a <=( A302  and  A299 );
 a21531a <=( (not A298)  and  a21530a );
 a21532a <=( a21531a  and  a21526a );
 a21535a <=( (not A169)  and  (not A170) );
 a21539a <=( A232  and  A202 );
 a21540a <=( (not A168)  and  a21539a );
 a21541a <=( a21540a  and  a21535a );
 a21544a <=( A236  and  (not A233) );
 a21548a <=( A269  and  A266 );
 a21549a <=( (not A265)  and  a21548a );
 a21550a <=( a21549a  and  a21544a );
 a21553a <=( (not A169)  and  (not A170) );
 a21557a <=( A232  and  A202 );
 a21558a <=( (not A168)  and  a21557a );
 a21559a <=( a21558a  and  a21553a );
 a21562a <=( A236  and  (not A233) );
 a21566a <=( A269  and  (not A266) );
 a21567a <=( A265  and  a21566a );
 a21568a <=( a21567a  and  a21562a );
 a21571a <=( (not A169)  and  (not A170) );
 a21575a <=( A201  and  A199 );
 a21576a <=( (not A168)  and  a21575a );
 a21577a <=( a21576a  and  a21571a );
 a21580a <=( A234  and  A232 );
 a21584a <=( A302  and  (not A299) );
 a21585a <=( A298  and  a21584a );
 a21586a <=( a21585a  and  a21580a );
 a21589a <=( (not A169)  and  (not A170) );
 a21593a <=( A201  and  A199 );
 a21594a <=( (not A168)  and  a21593a );
 a21595a <=( a21594a  and  a21589a );
 a21598a <=( A234  and  A232 );
 a21602a <=( A302  and  A299 );
 a21603a <=( (not A298)  and  a21602a );
 a21604a <=( a21603a  and  a21598a );
 a21607a <=( (not A169)  and  (not A170) );
 a21611a <=( A201  and  A199 );
 a21612a <=( (not A168)  and  a21611a );
 a21613a <=( a21612a  and  a21607a );
 a21616a <=( A234  and  A232 );
 a21620a <=( A269  and  A266 );
 a21621a <=( (not A265)  and  a21620a );
 a21622a <=( a21621a  and  a21616a );
 a21625a <=( (not A169)  and  (not A170) );
 a21629a <=( A201  and  A199 );
 a21630a <=( (not A168)  and  a21629a );
 a21631a <=( a21630a  and  a21625a );
 a21634a <=( A234  and  A232 );
 a21638a <=( A269  and  (not A266) );
 a21639a <=( A265  and  a21638a );
 a21640a <=( a21639a  and  a21634a );
 a21643a <=( (not A169)  and  (not A170) );
 a21647a <=( A201  and  A199 );
 a21648a <=( (not A168)  and  a21647a );
 a21649a <=( a21648a  and  a21643a );
 a21652a <=( A234  and  A233 );
 a21656a <=( A302  and  (not A299) );
 a21657a <=( A298  and  a21656a );
 a21658a <=( a21657a  and  a21652a );
 a21661a <=( (not A169)  and  (not A170) );
 a21665a <=( A201  and  A199 );
 a21666a <=( (not A168)  and  a21665a );
 a21667a <=( a21666a  and  a21661a );
 a21670a <=( A234  and  A233 );
 a21674a <=( A302  and  A299 );
 a21675a <=( (not A298)  and  a21674a );
 a21676a <=( a21675a  and  a21670a );
 a21679a <=( (not A169)  and  (not A170) );
 a21683a <=( A201  and  A199 );
 a21684a <=( (not A168)  and  a21683a );
 a21685a <=( a21684a  and  a21679a );
 a21688a <=( A234  and  A233 );
 a21692a <=( A269  and  A266 );
 a21693a <=( (not A265)  and  a21692a );
 a21694a <=( a21693a  and  a21688a );
 a21697a <=( (not A169)  and  (not A170) );
 a21701a <=( A201  and  A199 );
 a21702a <=( (not A168)  and  a21701a );
 a21703a <=( a21702a  and  a21697a );
 a21706a <=( A234  and  A233 );
 a21710a <=( A269  and  (not A266) );
 a21711a <=( A265  and  a21710a );
 a21712a <=( a21711a  and  a21706a );
 a21715a <=( (not A169)  and  (not A170) );
 a21719a <=( A201  and  A199 );
 a21720a <=( (not A168)  and  a21719a );
 a21721a <=( a21720a  and  a21715a );
 a21724a <=( A233  and  (not A232) );
 a21728a <=( A300  and  A299 );
 a21729a <=( A236  and  a21728a );
 a21730a <=( a21729a  and  a21724a );
 a21733a <=( (not A169)  and  (not A170) );
 a21737a <=( A201  and  A199 );
 a21738a <=( (not A168)  and  a21737a );
 a21739a <=( a21738a  and  a21733a );
 a21742a <=( A233  and  (not A232) );
 a21746a <=( A300  and  A298 );
 a21747a <=( A236  and  a21746a );
 a21748a <=( a21747a  and  a21742a );
 a21751a <=( (not A169)  and  (not A170) );
 a21755a <=( A201  and  A199 );
 a21756a <=( (not A168)  and  a21755a );
 a21757a <=( a21756a  and  a21751a );
 a21760a <=( A233  and  (not A232) );
 a21764a <=( A267  and  A265 );
 a21765a <=( A236  and  a21764a );
 a21766a <=( a21765a  and  a21760a );
 a21769a <=( (not A169)  and  (not A170) );
 a21773a <=( A201  and  A199 );
 a21774a <=( (not A168)  and  a21773a );
 a21775a <=( a21774a  and  a21769a );
 a21778a <=( A233  and  (not A232) );
 a21782a <=( A267  and  A266 );
 a21783a <=( A236  and  a21782a );
 a21784a <=( a21783a  and  a21778a );
 a21787a <=( (not A169)  and  (not A170) );
 a21791a <=( A201  and  A199 );
 a21792a <=( (not A168)  and  a21791a );
 a21793a <=( a21792a  and  a21787a );
 a21796a <=( (not A233)  and  A232 );
 a21800a <=( A300  and  A299 );
 a21801a <=( A236  and  a21800a );
 a21802a <=( a21801a  and  a21796a );
 a21805a <=( (not A169)  and  (not A170) );
 a21809a <=( A201  and  A199 );
 a21810a <=( (not A168)  and  a21809a );
 a21811a <=( a21810a  and  a21805a );
 a21814a <=( (not A233)  and  A232 );
 a21818a <=( A300  and  A298 );
 a21819a <=( A236  and  a21818a );
 a21820a <=( a21819a  and  a21814a );
 a21823a <=( (not A169)  and  (not A170) );
 a21827a <=( A201  and  A199 );
 a21828a <=( (not A168)  and  a21827a );
 a21829a <=( a21828a  and  a21823a );
 a21832a <=( (not A233)  and  A232 );
 a21836a <=( A267  and  A265 );
 a21837a <=( A236  and  a21836a );
 a21838a <=( a21837a  and  a21832a );
 a21841a <=( (not A169)  and  (not A170) );
 a21845a <=( A201  and  A199 );
 a21846a <=( (not A168)  and  a21845a );
 a21847a <=( a21846a  and  a21841a );
 a21850a <=( (not A233)  and  A232 );
 a21854a <=( A267  and  A266 );
 a21855a <=( A236  and  a21854a );
 a21856a <=( a21855a  and  a21850a );
 a21859a <=( (not A169)  and  (not A170) );
 a21863a <=( A201  and  A200 );
 a21864a <=( (not A168)  and  a21863a );
 a21865a <=( a21864a  and  a21859a );
 a21868a <=( A234  and  A232 );
 a21872a <=( A302  and  (not A299) );
 a21873a <=( A298  and  a21872a );
 a21874a <=( a21873a  and  a21868a );
 a21877a <=( (not A169)  and  (not A170) );
 a21881a <=( A201  and  A200 );
 a21882a <=( (not A168)  and  a21881a );
 a21883a <=( a21882a  and  a21877a );
 a21886a <=( A234  and  A232 );
 a21890a <=( A302  and  A299 );
 a21891a <=( (not A298)  and  a21890a );
 a21892a <=( a21891a  and  a21886a );
 a21895a <=( (not A169)  and  (not A170) );
 a21899a <=( A201  and  A200 );
 a21900a <=( (not A168)  and  a21899a );
 a21901a <=( a21900a  and  a21895a );
 a21904a <=( A234  and  A232 );
 a21908a <=( A269  and  A266 );
 a21909a <=( (not A265)  and  a21908a );
 a21910a <=( a21909a  and  a21904a );
 a21913a <=( (not A169)  and  (not A170) );
 a21917a <=( A201  and  A200 );
 a21918a <=( (not A168)  and  a21917a );
 a21919a <=( a21918a  and  a21913a );
 a21922a <=( A234  and  A232 );
 a21926a <=( A269  and  (not A266) );
 a21927a <=( A265  and  a21926a );
 a21928a <=( a21927a  and  a21922a );
 a21931a <=( (not A169)  and  (not A170) );
 a21935a <=( A201  and  A200 );
 a21936a <=( (not A168)  and  a21935a );
 a21937a <=( a21936a  and  a21931a );
 a21940a <=( A234  and  A233 );
 a21944a <=( A302  and  (not A299) );
 a21945a <=( A298  and  a21944a );
 a21946a <=( a21945a  and  a21940a );
 a21949a <=( (not A169)  and  (not A170) );
 a21953a <=( A201  and  A200 );
 a21954a <=( (not A168)  and  a21953a );
 a21955a <=( a21954a  and  a21949a );
 a21958a <=( A234  and  A233 );
 a21962a <=( A302  and  A299 );
 a21963a <=( (not A298)  and  a21962a );
 a21964a <=( a21963a  and  a21958a );
 a21967a <=( (not A169)  and  (not A170) );
 a21971a <=( A201  and  A200 );
 a21972a <=( (not A168)  and  a21971a );
 a21973a <=( a21972a  and  a21967a );
 a21976a <=( A234  and  A233 );
 a21980a <=( A269  and  A266 );
 a21981a <=( (not A265)  and  a21980a );
 a21982a <=( a21981a  and  a21976a );
 a21985a <=( (not A169)  and  (not A170) );
 a21989a <=( A201  and  A200 );
 a21990a <=( (not A168)  and  a21989a );
 a21991a <=( a21990a  and  a21985a );
 a21994a <=( A234  and  A233 );
 a21998a <=( A269  and  (not A266) );
 a21999a <=( A265  and  a21998a );
 a22000a <=( a21999a  and  a21994a );
 a22003a <=( (not A169)  and  (not A170) );
 a22007a <=( A201  and  A200 );
 a22008a <=( (not A168)  and  a22007a );
 a22009a <=( a22008a  and  a22003a );
 a22012a <=( A233  and  (not A232) );
 a22016a <=( A300  and  A299 );
 a22017a <=( A236  and  a22016a );
 a22018a <=( a22017a  and  a22012a );
 a22021a <=( (not A169)  and  (not A170) );
 a22025a <=( A201  and  A200 );
 a22026a <=( (not A168)  and  a22025a );
 a22027a <=( a22026a  and  a22021a );
 a22030a <=( A233  and  (not A232) );
 a22034a <=( A300  and  A298 );
 a22035a <=( A236  and  a22034a );
 a22036a <=( a22035a  and  a22030a );
 a22039a <=( (not A169)  and  (not A170) );
 a22043a <=( A201  and  A200 );
 a22044a <=( (not A168)  and  a22043a );
 a22045a <=( a22044a  and  a22039a );
 a22048a <=( A233  and  (not A232) );
 a22052a <=( A267  and  A265 );
 a22053a <=( A236  and  a22052a );
 a22054a <=( a22053a  and  a22048a );
 a22057a <=( (not A169)  and  (not A170) );
 a22061a <=( A201  and  A200 );
 a22062a <=( (not A168)  and  a22061a );
 a22063a <=( a22062a  and  a22057a );
 a22066a <=( A233  and  (not A232) );
 a22070a <=( A267  and  A266 );
 a22071a <=( A236  and  a22070a );
 a22072a <=( a22071a  and  a22066a );
 a22075a <=( (not A169)  and  (not A170) );
 a22079a <=( A201  and  A200 );
 a22080a <=( (not A168)  and  a22079a );
 a22081a <=( a22080a  and  a22075a );
 a22084a <=( (not A233)  and  A232 );
 a22088a <=( A300  and  A299 );
 a22089a <=( A236  and  a22088a );
 a22090a <=( a22089a  and  a22084a );
 a22093a <=( (not A169)  and  (not A170) );
 a22097a <=( A201  and  A200 );
 a22098a <=( (not A168)  and  a22097a );
 a22099a <=( a22098a  and  a22093a );
 a22102a <=( (not A233)  and  A232 );
 a22106a <=( A300  and  A298 );
 a22107a <=( A236  and  a22106a );
 a22108a <=( a22107a  and  a22102a );
 a22111a <=( (not A169)  and  (not A170) );
 a22115a <=( A201  and  A200 );
 a22116a <=( (not A168)  and  a22115a );
 a22117a <=( a22116a  and  a22111a );
 a22120a <=( (not A233)  and  A232 );
 a22124a <=( A267  and  A265 );
 a22125a <=( A236  and  a22124a );
 a22126a <=( a22125a  and  a22120a );
 a22129a <=( (not A169)  and  (not A170) );
 a22133a <=( A201  and  A200 );
 a22134a <=( (not A168)  and  a22133a );
 a22135a <=( a22134a  and  a22129a );
 a22138a <=( (not A233)  and  A232 );
 a22142a <=( A267  and  A266 );
 a22143a <=( A236  and  a22142a );
 a22144a <=( a22143a  and  a22138a );
 a22147a <=( (not A169)  and  (not A170) );
 a22151a <=( A200  and  (not A199) );
 a22152a <=( (not A168)  and  a22151a );
 a22153a <=( a22152a  and  a22147a );
 a22156a <=( A235  and  A203 );
 a22160a <=( A302  and  (not A299) );
 a22161a <=( A298  and  a22160a );
 a22162a <=( a22161a  and  a22156a );
 a22165a <=( (not A169)  and  (not A170) );
 a22169a <=( A200  and  (not A199) );
 a22170a <=( (not A168)  and  a22169a );
 a22171a <=( a22170a  and  a22165a );
 a22174a <=( A235  and  A203 );
 a22178a <=( A302  and  A299 );
 a22179a <=( (not A298)  and  a22178a );
 a22180a <=( a22179a  and  a22174a );
 a22183a <=( (not A169)  and  (not A170) );
 a22187a <=( A200  and  (not A199) );
 a22188a <=( (not A168)  and  a22187a );
 a22189a <=( a22188a  and  a22183a );
 a22192a <=( A235  and  A203 );
 a22196a <=( A269  and  A266 );
 a22197a <=( (not A265)  and  a22196a );
 a22198a <=( a22197a  and  a22192a );
 a22201a <=( (not A169)  and  (not A170) );
 a22205a <=( A200  and  (not A199) );
 a22206a <=( (not A168)  and  a22205a );
 a22207a <=( a22206a  and  a22201a );
 a22210a <=( A235  and  A203 );
 a22214a <=( A269  and  (not A266) );
 a22215a <=( A265  and  a22214a );
 a22216a <=( a22215a  and  a22210a );
 a22219a <=( (not A169)  and  (not A170) );
 a22223a <=( A200  and  (not A199) );
 a22224a <=( (not A168)  and  a22223a );
 a22225a <=( a22224a  and  a22219a );
 a22228a <=( A232  and  A203 );
 a22232a <=( A300  and  A299 );
 a22233a <=( A234  and  a22232a );
 a22234a <=( a22233a  and  a22228a );
 a22237a <=( (not A169)  and  (not A170) );
 a22241a <=( A200  and  (not A199) );
 a22242a <=( (not A168)  and  a22241a );
 a22243a <=( a22242a  and  a22237a );
 a22246a <=( A232  and  A203 );
 a22250a <=( A300  and  A298 );
 a22251a <=( A234  and  a22250a );
 a22252a <=( a22251a  and  a22246a );
 a22255a <=( (not A169)  and  (not A170) );
 a22259a <=( A200  and  (not A199) );
 a22260a <=( (not A168)  and  a22259a );
 a22261a <=( a22260a  and  a22255a );
 a22264a <=( A232  and  A203 );
 a22268a <=( A267  and  A265 );
 a22269a <=( A234  and  a22268a );
 a22270a <=( a22269a  and  a22264a );
 a22273a <=( (not A169)  and  (not A170) );
 a22277a <=( A200  and  (not A199) );
 a22278a <=( (not A168)  and  a22277a );
 a22279a <=( a22278a  and  a22273a );
 a22282a <=( A232  and  A203 );
 a22286a <=( A267  and  A266 );
 a22287a <=( A234  and  a22286a );
 a22288a <=( a22287a  and  a22282a );
 a22291a <=( (not A169)  and  (not A170) );
 a22295a <=( A200  and  (not A199) );
 a22296a <=( (not A168)  and  a22295a );
 a22297a <=( a22296a  and  a22291a );
 a22300a <=( A233  and  A203 );
 a22304a <=( A300  and  A299 );
 a22305a <=( A234  and  a22304a );
 a22306a <=( a22305a  and  a22300a );
 a22309a <=( (not A169)  and  (not A170) );
 a22313a <=( A200  and  (not A199) );
 a22314a <=( (not A168)  and  a22313a );
 a22315a <=( a22314a  and  a22309a );
 a22318a <=( A233  and  A203 );
 a22322a <=( A300  and  A298 );
 a22323a <=( A234  and  a22322a );
 a22324a <=( a22323a  and  a22318a );
 a22327a <=( (not A169)  and  (not A170) );
 a22331a <=( A200  and  (not A199) );
 a22332a <=( (not A168)  and  a22331a );
 a22333a <=( a22332a  and  a22327a );
 a22336a <=( A233  and  A203 );
 a22340a <=( A267  and  A265 );
 a22341a <=( A234  and  a22340a );
 a22342a <=( a22341a  and  a22336a );
 a22345a <=( (not A169)  and  (not A170) );
 a22349a <=( A200  and  (not A199) );
 a22350a <=( (not A168)  and  a22349a );
 a22351a <=( a22350a  and  a22345a );
 a22354a <=( A233  and  A203 );
 a22358a <=( A267  and  A266 );
 a22359a <=( A234  and  a22358a );
 a22360a <=( a22359a  and  a22354a );
 a22363a <=( (not A169)  and  (not A170) );
 a22367a <=( A200  and  (not A199) );
 a22368a <=( (not A168)  and  a22367a );
 a22369a <=( a22368a  and  a22363a );
 a22372a <=( (not A232)  and  A203 );
 a22376a <=( A301  and  A236 );
 a22377a <=( A233  and  a22376a );
 a22378a <=( a22377a  and  a22372a );
 a22381a <=( (not A169)  and  (not A170) );
 a22385a <=( A200  and  (not A199) );
 a22386a <=( (not A168)  and  a22385a );
 a22387a <=( a22386a  and  a22381a );
 a22390a <=( (not A232)  and  A203 );
 a22394a <=( A268  and  A236 );
 a22395a <=( A233  and  a22394a );
 a22396a <=( a22395a  and  a22390a );
 a22399a <=( (not A169)  and  (not A170) );
 a22403a <=( A200  and  (not A199) );
 a22404a <=( (not A168)  and  a22403a );
 a22405a <=( a22404a  and  a22399a );
 a22408a <=( A232  and  A203 );
 a22412a <=( A301  and  A236 );
 a22413a <=( (not A233)  and  a22412a );
 a22414a <=( a22413a  and  a22408a );
 a22417a <=( (not A169)  and  (not A170) );
 a22421a <=( A200  and  (not A199) );
 a22422a <=( (not A168)  and  a22421a );
 a22423a <=( a22422a  and  a22417a );
 a22426a <=( A232  and  A203 );
 a22430a <=( A268  and  A236 );
 a22431a <=( (not A233)  and  a22430a );
 a22432a <=( a22431a  and  a22426a );
 a22435a <=( (not A169)  and  (not A170) );
 a22439a <=( (not A200)  and  A199 );
 a22440a <=( (not A168)  and  a22439a );
 a22441a <=( a22440a  and  a22435a );
 a22444a <=( A235  and  A203 );
 a22448a <=( A302  and  (not A299) );
 a22449a <=( A298  and  a22448a );
 a22450a <=( a22449a  and  a22444a );
 a22453a <=( (not A169)  and  (not A170) );
 a22457a <=( (not A200)  and  A199 );
 a22458a <=( (not A168)  and  a22457a );
 a22459a <=( a22458a  and  a22453a );
 a22462a <=( A235  and  A203 );
 a22466a <=( A302  and  A299 );
 a22467a <=( (not A298)  and  a22466a );
 a22468a <=( a22467a  and  a22462a );
 a22471a <=( (not A169)  and  (not A170) );
 a22475a <=( (not A200)  and  A199 );
 a22476a <=( (not A168)  and  a22475a );
 a22477a <=( a22476a  and  a22471a );
 a22480a <=( A235  and  A203 );
 a22484a <=( A269  and  A266 );
 a22485a <=( (not A265)  and  a22484a );
 a22486a <=( a22485a  and  a22480a );
 a22489a <=( (not A169)  and  (not A170) );
 a22493a <=( (not A200)  and  A199 );
 a22494a <=( (not A168)  and  a22493a );
 a22495a <=( a22494a  and  a22489a );
 a22498a <=( A235  and  A203 );
 a22502a <=( A269  and  (not A266) );
 a22503a <=( A265  and  a22502a );
 a22504a <=( a22503a  and  a22498a );
 a22507a <=( (not A169)  and  (not A170) );
 a22511a <=( (not A200)  and  A199 );
 a22512a <=( (not A168)  and  a22511a );
 a22513a <=( a22512a  and  a22507a );
 a22516a <=( A232  and  A203 );
 a22520a <=( A300  and  A299 );
 a22521a <=( A234  and  a22520a );
 a22522a <=( a22521a  and  a22516a );
 a22525a <=( (not A169)  and  (not A170) );
 a22529a <=( (not A200)  and  A199 );
 a22530a <=( (not A168)  and  a22529a );
 a22531a <=( a22530a  and  a22525a );
 a22534a <=( A232  and  A203 );
 a22538a <=( A300  and  A298 );
 a22539a <=( A234  and  a22538a );
 a22540a <=( a22539a  and  a22534a );
 a22543a <=( (not A169)  and  (not A170) );
 a22547a <=( (not A200)  and  A199 );
 a22548a <=( (not A168)  and  a22547a );
 a22549a <=( a22548a  and  a22543a );
 a22552a <=( A232  and  A203 );
 a22556a <=( A267  and  A265 );
 a22557a <=( A234  and  a22556a );
 a22558a <=( a22557a  and  a22552a );
 a22561a <=( (not A169)  and  (not A170) );
 a22565a <=( (not A200)  and  A199 );
 a22566a <=( (not A168)  and  a22565a );
 a22567a <=( a22566a  and  a22561a );
 a22570a <=( A232  and  A203 );
 a22574a <=( A267  and  A266 );
 a22575a <=( A234  and  a22574a );
 a22576a <=( a22575a  and  a22570a );
 a22579a <=( (not A169)  and  (not A170) );
 a22583a <=( (not A200)  and  A199 );
 a22584a <=( (not A168)  and  a22583a );
 a22585a <=( a22584a  and  a22579a );
 a22588a <=( A233  and  A203 );
 a22592a <=( A300  and  A299 );
 a22593a <=( A234  and  a22592a );
 a22594a <=( a22593a  and  a22588a );
 a22597a <=( (not A169)  and  (not A170) );
 a22601a <=( (not A200)  and  A199 );
 a22602a <=( (not A168)  and  a22601a );
 a22603a <=( a22602a  and  a22597a );
 a22606a <=( A233  and  A203 );
 a22610a <=( A300  and  A298 );
 a22611a <=( A234  and  a22610a );
 a22612a <=( a22611a  and  a22606a );
 a22615a <=( (not A169)  and  (not A170) );
 a22619a <=( (not A200)  and  A199 );
 a22620a <=( (not A168)  and  a22619a );
 a22621a <=( a22620a  and  a22615a );
 a22624a <=( A233  and  A203 );
 a22628a <=( A267  and  A265 );
 a22629a <=( A234  and  a22628a );
 a22630a <=( a22629a  and  a22624a );
 a22633a <=( (not A169)  and  (not A170) );
 a22637a <=( (not A200)  and  A199 );
 a22638a <=( (not A168)  and  a22637a );
 a22639a <=( a22638a  and  a22633a );
 a22642a <=( A233  and  A203 );
 a22646a <=( A267  and  A266 );
 a22647a <=( A234  and  a22646a );
 a22648a <=( a22647a  and  a22642a );
 a22651a <=( (not A169)  and  (not A170) );
 a22655a <=( (not A200)  and  A199 );
 a22656a <=( (not A168)  and  a22655a );
 a22657a <=( a22656a  and  a22651a );
 a22660a <=( (not A232)  and  A203 );
 a22664a <=( A301  and  A236 );
 a22665a <=( A233  and  a22664a );
 a22666a <=( a22665a  and  a22660a );
 a22669a <=( (not A169)  and  (not A170) );
 a22673a <=( (not A200)  and  A199 );
 a22674a <=( (not A168)  and  a22673a );
 a22675a <=( a22674a  and  a22669a );
 a22678a <=( (not A232)  and  A203 );
 a22682a <=( A268  and  A236 );
 a22683a <=( A233  and  a22682a );
 a22684a <=( a22683a  and  a22678a );
 a22687a <=( (not A169)  and  (not A170) );
 a22691a <=( (not A200)  and  A199 );
 a22692a <=( (not A168)  and  a22691a );
 a22693a <=( a22692a  and  a22687a );
 a22696a <=( A232  and  A203 );
 a22700a <=( A301  and  A236 );
 a22701a <=( (not A233)  and  a22700a );
 a22702a <=( a22701a  and  a22696a );
 a22705a <=( (not A169)  and  (not A170) );
 a22709a <=( (not A200)  and  A199 );
 a22710a <=( (not A168)  and  a22709a );
 a22711a <=( a22710a  and  a22705a );
 a22714a <=( A232  and  A203 );
 a22718a <=( A268  and  A236 );
 a22719a <=( (not A233)  and  a22718a );
 a22720a <=( a22719a  and  a22714a );
 a22723a <=( A166  and  A168 );
 a22727a <=( (not A203)  and  (not A202) );
 a22728a <=( (not A201)  and  a22727a );
 a22729a <=( a22728a  and  a22723a );
 a22733a <=( A236  and  A233 );
 a22734a <=( (not A232)  and  a22733a );
 a22738a <=( A302  and  (not A299) );
 a22739a <=( A298  and  a22738a );
 a22740a <=( a22739a  and  a22734a );
 a22743a <=( A166  and  A168 );
 a22747a <=( (not A203)  and  (not A202) );
 a22748a <=( (not A201)  and  a22747a );
 a22749a <=( a22748a  and  a22743a );
 a22753a <=( A236  and  A233 );
 a22754a <=( (not A232)  and  a22753a );
 a22758a <=( A302  and  A299 );
 a22759a <=( (not A298)  and  a22758a );
 a22760a <=( a22759a  and  a22754a );
 a22763a <=( A166  and  A168 );
 a22767a <=( (not A203)  and  (not A202) );
 a22768a <=( (not A201)  and  a22767a );
 a22769a <=( a22768a  and  a22763a );
 a22773a <=( A236  and  A233 );
 a22774a <=( (not A232)  and  a22773a );
 a22778a <=( A269  and  A266 );
 a22779a <=( (not A265)  and  a22778a );
 a22780a <=( a22779a  and  a22774a );
 a22783a <=( A166  and  A168 );
 a22787a <=( (not A203)  and  (not A202) );
 a22788a <=( (not A201)  and  a22787a );
 a22789a <=( a22788a  and  a22783a );
 a22793a <=( A236  and  A233 );
 a22794a <=( (not A232)  and  a22793a );
 a22798a <=( A269  and  (not A266) );
 a22799a <=( A265  and  a22798a );
 a22800a <=( a22799a  and  a22794a );
 a22803a <=( A166  and  A168 );
 a22807a <=( (not A203)  and  (not A202) );
 a22808a <=( (not A201)  and  a22807a );
 a22809a <=( a22808a  and  a22803a );
 a22813a <=( A236  and  (not A233) );
 a22814a <=( A232  and  a22813a );
 a22818a <=( A302  and  (not A299) );
 a22819a <=( A298  and  a22818a );
 a22820a <=( a22819a  and  a22814a );
 a22823a <=( A166  and  A168 );
 a22827a <=( (not A203)  and  (not A202) );
 a22828a <=( (not A201)  and  a22827a );
 a22829a <=( a22828a  and  a22823a );
 a22833a <=( A236  and  (not A233) );
 a22834a <=( A232  and  a22833a );
 a22838a <=( A302  and  A299 );
 a22839a <=( (not A298)  and  a22838a );
 a22840a <=( a22839a  and  a22834a );
 a22843a <=( A166  and  A168 );
 a22847a <=( (not A203)  and  (not A202) );
 a22848a <=( (not A201)  and  a22847a );
 a22849a <=( a22848a  and  a22843a );
 a22853a <=( A236  and  (not A233) );
 a22854a <=( A232  and  a22853a );
 a22858a <=( A269  and  A266 );
 a22859a <=( (not A265)  and  a22858a );
 a22860a <=( a22859a  and  a22854a );
 a22863a <=( A166  and  A168 );
 a22867a <=( (not A203)  and  (not A202) );
 a22868a <=( (not A201)  and  a22867a );
 a22869a <=( a22868a  and  a22863a );
 a22873a <=( A236  and  (not A233) );
 a22874a <=( A232  and  a22873a );
 a22878a <=( A269  and  (not A266) );
 a22879a <=( A265  and  a22878a );
 a22880a <=( a22879a  and  a22874a );
 a22883a <=( A166  and  A168 );
 a22887a <=( (not A201)  and  A200 );
 a22888a <=( A199  and  a22887a );
 a22889a <=( a22888a  and  a22883a );
 a22893a <=( A234  and  A232 );
 a22894a <=( (not A202)  and  a22893a );
 a22898a <=( A302  and  (not A299) );
 a22899a <=( A298  and  a22898a );
 a22900a <=( a22899a  and  a22894a );
 a22903a <=( A166  and  A168 );
 a22907a <=( (not A201)  and  A200 );
 a22908a <=( A199  and  a22907a );
 a22909a <=( a22908a  and  a22903a );
 a22913a <=( A234  and  A232 );
 a22914a <=( (not A202)  and  a22913a );
 a22918a <=( A302  and  A299 );
 a22919a <=( (not A298)  and  a22918a );
 a22920a <=( a22919a  and  a22914a );
 a22923a <=( A166  and  A168 );
 a22927a <=( (not A201)  and  A200 );
 a22928a <=( A199  and  a22927a );
 a22929a <=( a22928a  and  a22923a );
 a22933a <=( A234  and  A232 );
 a22934a <=( (not A202)  and  a22933a );
 a22938a <=( A269  and  A266 );
 a22939a <=( (not A265)  and  a22938a );
 a22940a <=( a22939a  and  a22934a );
 a22943a <=( A166  and  A168 );
 a22947a <=( (not A201)  and  A200 );
 a22948a <=( A199  and  a22947a );
 a22949a <=( a22948a  and  a22943a );
 a22953a <=( A234  and  A232 );
 a22954a <=( (not A202)  and  a22953a );
 a22958a <=( A269  and  (not A266) );
 a22959a <=( A265  and  a22958a );
 a22960a <=( a22959a  and  a22954a );
 a22963a <=( A166  and  A168 );
 a22967a <=( (not A201)  and  A200 );
 a22968a <=( A199  and  a22967a );
 a22969a <=( a22968a  and  a22963a );
 a22973a <=( A234  and  A233 );
 a22974a <=( (not A202)  and  a22973a );
 a22978a <=( A302  and  (not A299) );
 a22979a <=( A298  and  a22978a );
 a22980a <=( a22979a  and  a22974a );
 a22983a <=( A166  and  A168 );
 a22987a <=( (not A201)  and  A200 );
 a22988a <=( A199  and  a22987a );
 a22989a <=( a22988a  and  a22983a );
 a22993a <=( A234  and  A233 );
 a22994a <=( (not A202)  and  a22993a );
 a22998a <=( A302  and  A299 );
 a22999a <=( (not A298)  and  a22998a );
 a23000a <=( a22999a  and  a22994a );
 a23003a <=( A166  and  A168 );
 a23007a <=( (not A201)  and  A200 );
 a23008a <=( A199  and  a23007a );
 a23009a <=( a23008a  and  a23003a );
 a23013a <=( A234  and  A233 );
 a23014a <=( (not A202)  and  a23013a );
 a23018a <=( A269  and  A266 );
 a23019a <=( (not A265)  and  a23018a );
 a23020a <=( a23019a  and  a23014a );
 a23023a <=( A166  and  A168 );
 a23027a <=( (not A201)  and  A200 );
 a23028a <=( A199  and  a23027a );
 a23029a <=( a23028a  and  a23023a );
 a23033a <=( A234  and  A233 );
 a23034a <=( (not A202)  and  a23033a );
 a23038a <=( A269  and  (not A266) );
 a23039a <=( A265  and  a23038a );
 a23040a <=( a23039a  and  a23034a );
 a23043a <=( A166  and  A168 );
 a23047a <=( (not A201)  and  A200 );
 a23048a <=( A199  and  a23047a );
 a23049a <=( a23048a  and  a23043a );
 a23053a <=( A233  and  (not A232) );
 a23054a <=( (not A202)  and  a23053a );
 a23058a <=( A300  and  A299 );
 a23059a <=( A236  and  a23058a );
 a23060a <=( a23059a  and  a23054a );
 a23063a <=( A166  and  A168 );
 a23067a <=( (not A201)  and  A200 );
 a23068a <=( A199  and  a23067a );
 a23069a <=( a23068a  and  a23063a );
 a23073a <=( A233  and  (not A232) );
 a23074a <=( (not A202)  and  a23073a );
 a23078a <=( A300  and  A298 );
 a23079a <=( A236  and  a23078a );
 a23080a <=( a23079a  and  a23074a );
 a23083a <=( A166  and  A168 );
 a23087a <=( (not A201)  and  A200 );
 a23088a <=( A199  and  a23087a );
 a23089a <=( a23088a  and  a23083a );
 a23093a <=( A233  and  (not A232) );
 a23094a <=( (not A202)  and  a23093a );
 a23098a <=( A267  and  A265 );
 a23099a <=( A236  and  a23098a );
 a23100a <=( a23099a  and  a23094a );
 a23103a <=( A166  and  A168 );
 a23107a <=( (not A201)  and  A200 );
 a23108a <=( A199  and  a23107a );
 a23109a <=( a23108a  and  a23103a );
 a23113a <=( A233  and  (not A232) );
 a23114a <=( (not A202)  and  a23113a );
 a23118a <=( A267  and  A266 );
 a23119a <=( A236  and  a23118a );
 a23120a <=( a23119a  and  a23114a );
 a23123a <=( A166  and  A168 );
 a23127a <=( (not A201)  and  A200 );
 a23128a <=( A199  and  a23127a );
 a23129a <=( a23128a  and  a23123a );
 a23133a <=( (not A233)  and  A232 );
 a23134a <=( (not A202)  and  a23133a );
 a23138a <=( A300  and  A299 );
 a23139a <=( A236  and  a23138a );
 a23140a <=( a23139a  and  a23134a );
 a23143a <=( A166  and  A168 );
 a23147a <=( (not A201)  and  A200 );
 a23148a <=( A199  and  a23147a );
 a23149a <=( a23148a  and  a23143a );
 a23153a <=( (not A233)  and  A232 );
 a23154a <=( (not A202)  and  a23153a );
 a23158a <=( A300  and  A298 );
 a23159a <=( A236  and  a23158a );
 a23160a <=( a23159a  and  a23154a );
 a23163a <=( A166  and  A168 );
 a23167a <=( (not A201)  and  A200 );
 a23168a <=( A199  and  a23167a );
 a23169a <=( a23168a  and  a23163a );
 a23173a <=( (not A233)  and  A232 );
 a23174a <=( (not A202)  and  a23173a );
 a23178a <=( A267  and  A265 );
 a23179a <=( A236  and  a23178a );
 a23180a <=( a23179a  and  a23174a );
 a23183a <=( A166  and  A168 );
 a23187a <=( (not A201)  and  A200 );
 a23188a <=( A199  and  a23187a );
 a23189a <=( a23188a  and  a23183a );
 a23193a <=( (not A233)  and  A232 );
 a23194a <=( (not A202)  and  a23193a );
 a23198a <=( A267  and  A266 );
 a23199a <=( A236  and  a23198a );
 a23200a <=( a23199a  and  a23194a );
 a23203a <=( A166  and  A168 );
 a23207a <=( (not A202)  and  (not A200) );
 a23208a <=( (not A199)  and  a23207a );
 a23209a <=( a23208a  and  a23203a );
 a23213a <=( A236  and  A233 );
 a23214a <=( (not A232)  and  a23213a );
 a23218a <=( A302  and  (not A299) );
 a23219a <=( A298  and  a23218a );
 a23220a <=( a23219a  and  a23214a );
 a23223a <=( A166  and  A168 );
 a23227a <=( (not A202)  and  (not A200) );
 a23228a <=( (not A199)  and  a23227a );
 a23229a <=( a23228a  and  a23223a );
 a23233a <=( A236  and  A233 );
 a23234a <=( (not A232)  and  a23233a );
 a23238a <=( A302  and  A299 );
 a23239a <=( (not A298)  and  a23238a );
 a23240a <=( a23239a  and  a23234a );
 a23243a <=( A166  and  A168 );
 a23247a <=( (not A202)  and  (not A200) );
 a23248a <=( (not A199)  and  a23247a );
 a23249a <=( a23248a  and  a23243a );
 a23253a <=( A236  and  A233 );
 a23254a <=( (not A232)  and  a23253a );
 a23258a <=( A269  and  A266 );
 a23259a <=( (not A265)  and  a23258a );
 a23260a <=( a23259a  and  a23254a );
 a23263a <=( A166  and  A168 );
 a23267a <=( (not A202)  and  (not A200) );
 a23268a <=( (not A199)  and  a23267a );
 a23269a <=( a23268a  and  a23263a );
 a23273a <=( A236  and  A233 );
 a23274a <=( (not A232)  and  a23273a );
 a23278a <=( A269  and  (not A266) );
 a23279a <=( A265  and  a23278a );
 a23280a <=( a23279a  and  a23274a );
 a23283a <=( A166  and  A168 );
 a23287a <=( (not A202)  and  (not A200) );
 a23288a <=( (not A199)  and  a23287a );
 a23289a <=( a23288a  and  a23283a );
 a23293a <=( A236  and  (not A233) );
 a23294a <=( A232  and  a23293a );
 a23298a <=( A302  and  (not A299) );
 a23299a <=( A298  and  a23298a );
 a23300a <=( a23299a  and  a23294a );
 a23303a <=( A166  and  A168 );
 a23307a <=( (not A202)  and  (not A200) );
 a23308a <=( (not A199)  and  a23307a );
 a23309a <=( a23308a  and  a23303a );
 a23313a <=( A236  and  (not A233) );
 a23314a <=( A232  and  a23313a );
 a23318a <=( A302  and  A299 );
 a23319a <=( (not A298)  and  a23318a );
 a23320a <=( a23319a  and  a23314a );
 a23323a <=( A166  and  A168 );
 a23327a <=( (not A202)  and  (not A200) );
 a23328a <=( (not A199)  and  a23327a );
 a23329a <=( a23328a  and  a23323a );
 a23333a <=( A236  and  (not A233) );
 a23334a <=( A232  and  a23333a );
 a23338a <=( A269  and  A266 );
 a23339a <=( (not A265)  and  a23338a );
 a23340a <=( a23339a  and  a23334a );
 a23343a <=( A166  and  A168 );
 a23347a <=( (not A202)  and  (not A200) );
 a23348a <=( (not A199)  and  a23347a );
 a23349a <=( a23348a  and  a23343a );
 a23353a <=( A236  and  (not A233) );
 a23354a <=( A232  and  a23353a );
 a23358a <=( A269  and  (not A266) );
 a23359a <=( A265  and  a23358a );
 a23360a <=( a23359a  and  a23354a );
 a23363a <=( A167  and  A168 );
 a23367a <=( (not A203)  and  (not A202) );
 a23368a <=( (not A201)  and  a23367a );
 a23369a <=( a23368a  and  a23363a );
 a23373a <=( A236  and  A233 );
 a23374a <=( (not A232)  and  a23373a );
 a23378a <=( A302  and  (not A299) );
 a23379a <=( A298  and  a23378a );
 a23380a <=( a23379a  and  a23374a );
 a23383a <=( A167  and  A168 );
 a23387a <=( (not A203)  and  (not A202) );
 a23388a <=( (not A201)  and  a23387a );
 a23389a <=( a23388a  and  a23383a );
 a23393a <=( A236  and  A233 );
 a23394a <=( (not A232)  and  a23393a );
 a23398a <=( A302  and  A299 );
 a23399a <=( (not A298)  and  a23398a );
 a23400a <=( a23399a  and  a23394a );
 a23403a <=( A167  and  A168 );
 a23407a <=( (not A203)  and  (not A202) );
 a23408a <=( (not A201)  and  a23407a );
 a23409a <=( a23408a  and  a23403a );
 a23413a <=( A236  and  A233 );
 a23414a <=( (not A232)  and  a23413a );
 a23418a <=( A269  and  A266 );
 a23419a <=( (not A265)  and  a23418a );
 a23420a <=( a23419a  and  a23414a );
 a23423a <=( A167  and  A168 );
 a23427a <=( (not A203)  and  (not A202) );
 a23428a <=( (not A201)  and  a23427a );
 a23429a <=( a23428a  and  a23423a );
 a23433a <=( A236  and  A233 );
 a23434a <=( (not A232)  and  a23433a );
 a23438a <=( A269  and  (not A266) );
 a23439a <=( A265  and  a23438a );
 a23440a <=( a23439a  and  a23434a );
 a23443a <=( A167  and  A168 );
 a23447a <=( (not A203)  and  (not A202) );
 a23448a <=( (not A201)  and  a23447a );
 a23449a <=( a23448a  and  a23443a );
 a23453a <=( A236  and  (not A233) );
 a23454a <=( A232  and  a23453a );
 a23458a <=( A302  and  (not A299) );
 a23459a <=( A298  and  a23458a );
 a23460a <=( a23459a  and  a23454a );
 a23463a <=( A167  and  A168 );
 a23467a <=( (not A203)  and  (not A202) );
 a23468a <=( (not A201)  and  a23467a );
 a23469a <=( a23468a  and  a23463a );
 a23473a <=( A236  and  (not A233) );
 a23474a <=( A232  and  a23473a );
 a23478a <=( A302  and  A299 );
 a23479a <=( (not A298)  and  a23478a );
 a23480a <=( a23479a  and  a23474a );
 a23483a <=( A167  and  A168 );
 a23487a <=( (not A203)  and  (not A202) );
 a23488a <=( (not A201)  and  a23487a );
 a23489a <=( a23488a  and  a23483a );
 a23493a <=( A236  and  (not A233) );
 a23494a <=( A232  and  a23493a );
 a23498a <=( A269  and  A266 );
 a23499a <=( (not A265)  and  a23498a );
 a23500a <=( a23499a  and  a23494a );
 a23503a <=( A167  and  A168 );
 a23507a <=( (not A203)  and  (not A202) );
 a23508a <=( (not A201)  and  a23507a );
 a23509a <=( a23508a  and  a23503a );
 a23513a <=( A236  and  (not A233) );
 a23514a <=( A232  and  a23513a );
 a23518a <=( A269  and  (not A266) );
 a23519a <=( A265  and  a23518a );
 a23520a <=( a23519a  and  a23514a );
 a23523a <=( A167  and  A168 );
 a23527a <=( (not A201)  and  A200 );
 a23528a <=( A199  and  a23527a );
 a23529a <=( a23528a  and  a23523a );
 a23533a <=( A234  and  A232 );
 a23534a <=( (not A202)  and  a23533a );
 a23538a <=( A302  and  (not A299) );
 a23539a <=( A298  and  a23538a );
 a23540a <=( a23539a  and  a23534a );
 a23543a <=( A167  and  A168 );
 a23547a <=( (not A201)  and  A200 );
 a23548a <=( A199  and  a23547a );
 a23549a <=( a23548a  and  a23543a );
 a23553a <=( A234  and  A232 );
 a23554a <=( (not A202)  and  a23553a );
 a23558a <=( A302  and  A299 );
 a23559a <=( (not A298)  and  a23558a );
 a23560a <=( a23559a  and  a23554a );
 a23563a <=( A167  and  A168 );
 a23567a <=( (not A201)  and  A200 );
 a23568a <=( A199  and  a23567a );
 a23569a <=( a23568a  and  a23563a );
 a23573a <=( A234  and  A232 );
 a23574a <=( (not A202)  and  a23573a );
 a23578a <=( A269  and  A266 );
 a23579a <=( (not A265)  and  a23578a );
 a23580a <=( a23579a  and  a23574a );
 a23583a <=( A167  and  A168 );
 a23587a <=( (not A201)  and  A200 );
 a23588a <=( A199  and  a23587a );
 a23589a <=( a23588a  and  a23583a );
 a23593a <=( A234  and  A232 );
 a23594a <=( (not A202)  and  a23593a );
 a23598a <=( A269  and  (not A266) );
 a23599a <=( A265  and  a23598a );
 a23600a <=( a23599a  and  a23594a );
 a23603a <=( A167  and  A168 );
 a23607a <=( (not A201)  and  A200 );
 a23608a <=( A199  and  a23607a );
 a23609a <=( a23608a  and  a23603a );
 a23613a <=( A234  and  A233 );
 a23614a <=( (not A202)  and  a23613a );
 a23618a <=( A302  and  (not A299) );
 a23619a <=( A298  and  a23618a );
 a23620a <=( a23619a  and  a23614a );
 a23623a <=( A167  and  A168 );
 a23627a <=( (not A201)  and  A200 );
 a23628a <=( A199  and  a23627a );
 a23629a <=( a23628a  and  a23623a );
 a23633a <=( A234  and  A233 );
 a23634a <=( (not A202)  and  a23633a );
 a23638a <=( A302  and  A299 );
 a23639a <=( (not A298)  and  a23638a );
 a23640a <=( a23639a  and  a23634a );
 a23643a <=( A167  and  A168 );
 a23647a <=( (not A201)  and  A200 );
 a23648a <=( A199  and  a23647a );
 a23649a <=( a23648a  and  a23643a );
 a23653a <=( A234  and  A233 );
 a23654a <=( (not A202)  and  a23653a );
 a23658a <=( A269  and  A266 );
 a23659a <=( (not A265)  and  a23658a );
 a23660a <=( a23659a  and  a23654a );
 a23663a <=( A167  and  A168 );
 a23667a <=( (not A201)  and  A200 );
 a23668a <=( A199  and  a23667a );
 a23669a <=( a23668a  and  a23663a );
 a23673a <=( A234  and  A233 );
 a23674a <=( (not A202)  and  a23673a );
 a23678a <=( A269  and  (not A266) );
 a23679a <=( A265  and  a23678a );
 a23680a <=( a23679a  and  a23674a );
 a23683a <=( A167  and  A168 );
 a23687a <=( (not A201)  and  A200 );
 a23688a <=( A199  and  a23687a );
 a23689a <=( a23688a  and  a23683a );
 a23693a <=( A233  and  (not A232) );
 a23694a <=( (not A202)  and  a23693a );
 a23698a <=( A300  and  A299 );
 a23699a <=( A236  and  a23698a );
 a23700a <=( a23699a  and  a23694a );
 a23703a <=( A167  and  A168 );
 a23707a <=( (not A201)  and  A200 );
 a23708a <=( A199  and  a23707a );
 a23709a <=( a23708a  and  a23703a );
 a23713a <=( A233  and  (not A232) );
 a23714a <=( (not A202)  and  a23713a );
 a23718a <=( A300  and  A298 );
 a23719a <=( A236  and  a23718a );
 a23720a <=( a23719a  and  a23714a );
 a23723a <=( A167  and  A168 );
 a23727a <=( (not A201)  and  A200 );
 a23728a <=( A199  and  a23727a );
 a23729a <=( a23728a  and  a23723a );
 a23733a <=( A233  and  (not A232) );
 a23734a <=( (not A202)  and  a23733a );
 a23738a <=( A267  and  A265 );
 a23739a <=( A236  and  a23738a );
 a23740a <=( a23739a  and  a23734a );
 a23743a <=( A167  and  A168 );
 a23747a <=( (not A201)  and  A200 );
 a23748a <=( A199  and  a23747a );
 a23749a <=( a23748a  and  a23743a );
 a23753a <=( A233  and  (not A232) );
 a23754a <=( (not A202)  and  a23753a );
 a23758a <=( A267  and  A266 );
 a23759a <=( A236  and  a23758a );
 a23760a <=( a23759a  and  a23754a );
 a23763a <=( A167  and  A168 );
 a23767a <=( (not A201)  and  A200 );
 a23768a <=( A199  and  a23767a );
 a23769a <=( a23768a  and  a23763a );
 a23773a <=( (not A233)  and  A232 );
 a23774a <=( (not A202)  and  a23773a );
 a23778a <=( A300  and  A299 );
 a23779a <=( A236  and  a23778a );
 a23780a <=( a23779a  and  a23774a );
 a23783a <=( A167  and  A168 );
 a23787a <=( (not A201)  and  A200 );
 a23788a <=( A199  and  a23787a );
 a23789a <=( a23788a  and  a23783a );
 a23793a <=( (not A233)  and  A232 );
 a23794a <=( (not A202)  and  a23793a );
 a23798a <=( A300  and  A298 );
 a23799a <=( A236  and  a23798a );
 a23800a <=( a23799a  and  a23794a );
 a23803a <=( A167  and  A168 );
 a23807a <=( (not A201)  and  A200 );
 a23808a <=( A199  and  a23807a );
 a23809a <=( a23808a  and  a23803a );
 a23813a <=( (not A233)  and  A232 );
 a23814a <=( (not A202)  and  a23813a );
 a23818a <=( A267  and  A265 );
 a23819a <=( A236  and  a23818a );
 a23820a <=( a23819a  and  a23814a );
 a23823a <=( A167  and  A168 );
 a23827a <=( (not A201)  and  A200 );
 a23828a <=( A199  and  a23827a );
 a23829a <=( a23828a  and  a23823a );
 a23833a <=( (not A233)  and  A232 );
 a23834a <=( (not A202)  and  a23833a );
 a23838a <=( A267  and  A266 );
 a23839a <=( A236  and  a23838a );
 a23840a <=( a23839a  and  a23834a );
 a23843a <=( A167  and  A168 );
 a23847a <=( (not A202)  and  (not A200) );
 a23848a <=( (not A199)  and  a23847a );
 a23849a <=( a23848a  and  a23843a );
 a23853a <=( A236  and  A233 );
 a23854a <=( (not A232)  and  a23853a );
 a23858a <=( A302  and  (not A299) );
 a23859a <=( A298  and  a23858a );
 a23860a <=( a23859a  and  a23854a );
 a23863a <=( A167  and  A168 );
 a23867a <=( (not A202)  and  (not A200) );
 a23868a <=( (not A199)  and  a23867a );
 a23869a <=( a23868a  and  a23863a );
 a23873a <=( A236  and  A233 );
 a23874a <=( (not A232)  and  a23873a );
 a23878a <=( A302  and  A299 );
 a23879a <=( (not A298)  and  a23878a );
 a23880a <=( a23879a  and  a23874a );
 a23883a <=( A167  and  A168 );
 a23887a <=( (not A202)  and  (not A200) );
 a23888a <=( (not A199)  and  a23887a );
 a23889a <=( a23888a  and  a23883a );
 a23893a <=( A236  and  A233 );
 a23894a <=( (not A232)  and  a23893a );
 a23898a <=( A269  and  A266 );
 a23899a <=( (not A265)  and  a23898a );
 a23900a <=( a23899a  and  a23894a );
 a23903a <=( A167  and  A168 );
 a23907a <=( (not A202)  and  (not A200) );
 a23908a <=( (not A199)  and  a23907a );
 a23909a <=( a23908a  and  a23903a );
 a23913a <=( A236  and  A233 );
 a23914a <=( (not A232)  and  a23913a );
 a23918a <=( A269  and  (not A266) );
 a23919a <=( A265  and  a23918a );
 a23920a <=( a23919a  and  a23914a );
 a23923a <=( A167  and  A168 );
 a23927a <=( (not A202)  and  (not A200) );
 a23928a <=( (not A199)  and  a23927a );
 a23929a <=( a23928a  and  a23923a );
 a23933a <=( A236  and  (not A233) );
 a23934a <=( A232  and  a23933a );
 a23938a <=( A302  and  (not A299) );
 a23939a <=( A298  and  a23938a );
 a23940a <=( a23939a  and  a23934a );
 a23943a <=( A167  and  A168 );
 a23947a <=( (not A202)  and  (not A200) );
 a23948a <=( (not A199)  and  a23947a );
 a23949a <=( a23948a  and  a23943a );
 a23953a <=( A236  and  (not A233) );
 a23954a <=( A232  and  a23953a );
 a23958a <=( A302  and  A299 );
 a23959a <=( (not A298)  and  a23958a );
 a23960a <=( a23959a  and  a23954a );
 a23963a <=( A167  and  A168 );
 a23967a <=( (not A202)  and  (not A200) );
 a23968a <=( (not A199)  and  a23967a );
 a23969a <=( a23968a  and  a23963a );
 a23973a <=( A236  and  (not A233) );
 a23974a <=( A232  and  a23973a );
 a23978a <=( A269  and  A266 );
 a23979a <=( (not A265)  and  a23978a );
 a23980a <=( a23979a  and  a23974a );
 a23983a <=( A167  and  A168 );
 a23987a <=( (not A202)  and  (not A200) );
 a23988a <=( (not A199)  and  a23987a );
 a23989a <=( a23988a  and  a23983a );
 a23993a <=( A236  and  (not A233) );
 a23994a <=( A232  and  a23993a );
 a23998a <=( A269  and  (not A266) );
 a23999a <=( A265  and  a23998a );
 a24000a <=( a23999a  and  a23994a );
 a24003a <=( A167  and  A170 );
 a24007a <=( (not A202)  and  (not A201) );
 a24008a <=( (not A166)  and  a24007a );
 a24009a <=( a24008a  and  a24003a );
 a24013a <=( A234  and  A232 );
 a24014a <=( (not A203)  and  a24013a );
 a24018a <=( A302  and  (not A299) );
 a24019a <=( A298  and  a24018a );
 a24020a <=( a24019a  and  a24014a );
 a24023a <=( A167  and  A170 );
 a24027a <=( (not A202)  and  (not A201) );
 a24028a <=( (not A166)  and  a24027a );
 a24029a <=( a24028a  and  a24023a );
 a24033a <=( A234  and  A232 );
 a24034a <=( (not A203)  and  a24033a );
 a24038a <=( A302  and  A299 );
 a24039a <=( (not A298)  and  a24038a );
 a24040a <=( a24039a  and  a24034a );
 a24043a <=( A167  and  A170 );
 a24047a <=( (not A202)  and  (not A201) );
 a24048a <=( (not A166)  and  a24047a );
 a24049a <=( a24048a  and  a24043a );
 a24053a <=( A234  and  A232 );
 a24054a <=( (not A203)  and  a24053a );
 a24058a <=( A269  and  A266 );
 a24059a <=( (not A265)  and  a24058a );
 a24060a <=( a24059a  and  a24054a );
 a24063a <=( A167  and  A170 );
 a24067a <=( (not A202)  and  (not A201) );
 a24068a <=( (not A166)  and  a24067a );
 a24069a <=( a24068a  and  a24063a );
 a24073a <=( A234  and  A232 );
 a24074a <=( (not A203)  and  a24073a );
 a24078a <=( A269  and  (not A266) );
 a24079a <=( A265  and  a24078a );
 a24080a <=( a24079a  and  a24074a );
 a24083a <=( A167  and  A170 );
 a24087a <=( (not A202)  and  (not A201) );
 a24088a <=( (not A166)  and  a24087a );
 a24089a <=( a24088a  and  a24083a );
 a24093a <=( A234  and  A233 );
 a24094a <=( (not A203)  and  a24093a );
 a24098a <=( A302  and  (not A299) );
 a24099a <=( A298  and  a24098a );
 a24100a <=( a24099a  and  a24094a );
 a24103a <=( A167  and  A170 );
 a24107a <=( (not A202)  and  (not A201) );
 a24108a <=( (not A166)  and  a24107a );
 a24109a <=( a24108a  and  a24103a );
 a24113a <=( A234  and  A233 );
 a24114a <=( (not A203)  and  a24113a );
 a24118a <=( A302  and  A299 );
 a24119a <=( (not A298)  and  a24118a );
 a24120a <=( a24119a  and  a24114a );
 a24123a <=( A167  and  A170 );
 a24127a <=( (not A202)  and  (not A201) );
 a24128a <=( (not A166)  and  a24127a );
 a24129a <=( a24128a  and  a24123a );
 a24133a <=( A234  and  A233 );
 a24134a <=( (not A203)  and  a24133a );
 a24138a <=( A269  and  A266 );
 a24139a <=( (not A265)  and  a24138a );
 a24140a <=( a24139a  and  a24134a );
 a24143a <=( A167  and  A170 );
 a24147a <=( (not A202)  and  (not A201) );
 a24148a <=( (not A166)  and  a24147a );
 a24149a <=( a24148a  and  a24143a );
 a24153a <=( A234  and  A233 );
 a24154a <=( (not A203)  and  a24153a );
 a24158a <=( A269  and  (not A266) );
 a24159a <=( A265  and  a24158a );
 a24160a <=( a24159a  and  a24154a );
 a24163a <=( A167  and  A170 );
 a24167a <=( (not A202)  and  (not A201) );
 a24168a <=( (not A166)  and  a24167a );
 a24169a <=( a24168a  and  a24163a );
 a24173a <=( A233  and  (not A232) );
 a24174a <=( (not A203)  and  a24173a );
 a24178a <=( A300  and  A299 );
 a24179a <=( A236  and  a24178a );
 a24180a <=( a24179a  and  a24174a );
 a24183a <=( A167  and  A170 );
 a24187a <=( (not A202)  and  (not A201) );
 a24188a <=( (not A166)  and  a24187a );
 a24189a <=( a24188a  and  a24183a );
 a24193a <=( A233  and  (not A232) );
 a24194a <=( (not A203)  and  a24193a );
 a24198a <=( A300  and  A298 );
 a24199a <=( A236  and  a24198a );
 a24200a <=( a24199a  and  a24194a );
 a24203a <=( A167  and  A170 );
 a24207a <=( (not A202)  and  (not A201) );
 a24208a <=( (not A166)  and  a24207a );
 a24209a <=( a24208a  and  a24203a );
 a24213a <=( A233  and  (not A232) );
 a24214a <=( (not A203)  and  a24213a );
 a24218a <=( A267  and  A265 );
 a24219a <=( A236  and  a24218a );
 a24220a <=( a24219a  and  a24214a );
 a24223a <=( A167  and  A170 );
 a24227a <=( (not A202)  and  (not A201) );
 a24228a <=( (not A166)  and  a24227a );
 a24229a <=( a24228a  and  a24223a );
 a24233a <=( A233  and  (not A232) );
 a24234a <=( (not A203)  and  a24233a );
 a24238a <=( A267  and  A266 );
 a24239a <=( A236  and  a24238a );
 a24240a <=( a24239a  and  a24234a );
 a24243a <=( A167  and  A170 );
 a24247a <=( (not A202)  and  (not A201) );
 a24248a <=( (not A166)  and  a24247a );
 a24249a <=( a24248a  and  a24243a );
 a24253a <=( (not A233)  and  A232 );
 a24254a <=( (not A203)  and  a24253a );
 a24258a <=( A300  and  A299 );
 a24259a <=( A236  and  a24258a );
 a24260a <=( a24259a  and  a24254a );
 a24263a <=( A167  and  A170 );
 a24267a <=( (not A202)  and  (not A201) );
 a24268a <=( (not A166)  and  a24267a );
 a24269a <=( a24268a  and  a24263a );
 a24273a <=( (not A233)  and  A232 );
 a24274a <=( (not A203)  and  a24273a );
 a24278a <=( A300  and  A298 );
 a24279a <=( A236  and  a24278a );
 a24280a <=( a24279a  and  a24274a );
 a24283a <=( A167  and  A170 );
 a24287a <=( (not A202)  and  (not A201) );
 a24288a <=( (not A166)  and  a24287a );
 a24289a <=( a24288a  and  a24283a );
 a24293a <=( (not A233)  and  A232 );
 a24294a <=( (not A203)  and  a24293a );
 a24298a <=( A267  and  A265 );
 a24299a <=( A236  and  a24298a );
 a24300a <=( a24299a  and  a24294a );
 a24303a <=( A167  and  A170 );
 a24307a <=( (not A202)  and  (not A201) );
 a24308a <=( (not A166)  and  a24307a );
 a24309a <=( a24308a  and  a24303a );
 a24313a <=( (not A233)  and  A232 );
 a24314a <=( (not A203)  and  a24313a );
 a24318a <=( A267  and  A266 );
 a24319a <=( A236  and  a24318a );
 a24320a <=( a24319a  and  a24314a );
 a24323a <=( A167  and  A170 );
 a24327a <=( A200  and  A199 );
 a24328a <=( (not A166)  and  a24327a );
 a24329a <=( a24328a  and  a24323a );
 a24333a <=( A235  and  (not A202) );
 a24334a <=( (not A201)  and  a24333a );
 a24338a <=( A302  and  (not A299) );
 a24339a <=( A298  and  a24338a );
 a24340a <=( a24339a  and  a24334a );
 a24343a <=( A167  and  A170 );
 a24347a <=( A200  and  A199 );
 a24348a <=( (not A166)  and  a24347a );
 a24349a <=( a24348a  and  a24343a );
 a24353a <=( A235  and  (not A202) );
 a24354a <=( (not A201)  and  a24353a );
 a24358a <=( A302  and  A299 );
 a24359a <=( (not A298)  and  a24358a );
 a24360a <=( a24359a  and  a24354a );
 a24363a <=( A167  and  A170 );
 a24367a <=( A200  and  A199 );
 a24368a <=( (not A166)  and  a24367a );
 a24369a <=( a24368a  and  a24363a );
 a24373a <=( A235  and  (not A202) );
 a24374a <=( (not A201)  and  a24373a );
 a24378a <=( A269  and  A266 );
 a24379a <=( (not A265)  and  a24378a );
 a24380a <=( a24379a  and  a24374a );
 a24383a <=( A167  and  A170 );
 a24387a <=( A200  and  A199 );
 a24388a <=( (not A166)  and  a24387a );
 a24389a <=( a24388a  and  a24383a );
 a24393a <=( A235  and  (not A202) );
 a24394a <=( (not A201)  and  a24393a );
 a24398a <=( A269  and  (not A266) );
 a24399a <=( A265  and  a24398a );
 a24400a <=( a24399a  and  a24394a );
 a24403a <=( A167  and  A170 );
 a24407a <=( A200  and  A199 );
 a24408a <=( (not A166)  and  a24407a );
 a24409a <=( a24408a  and  a24403a );
 a24413a <=( A232  and  (not A202) );
 a24414a <=( (not A201)  and  a24413a );
 a24418a <=( A300  and  A299 );
 a24419a <=( A234  and  a24418a );
 a24420a <=( a24419a  and  a24414a );
 a24423a <=( A167  and  A170 );
 a24427a <=( A200  and  A199 );
 a24428a <=( (not A166)  and  a24427a );
 a24429a <=( a24428a  and  a24423a );
 a24433a <=( A232  and  (not A202) );
 a24434a <=( (not A201)  and  a24433a );
 a24438a <=( A300  and  A298 );
 a24439a <=( A234  and  a24438a );
 a24440a <=( a24439a  and  a24434a );
 a24443a <=( A167  and  A170 );
 a24447a <=( A200  and  A199 );
 a24448a <=( (not A166)  and  a24447a );
 a24449a <=( a24448a  and  a24443a );
 a24453a <=( A232  and  (not A202) );
 a24454a <=( (not A201)  and  a24453a );
 a24458a <=( A267  and  A265 );
 a24459a <=( A234  and  a24458a );
 a24460a <=( a24459a  and  a24454a );
 a24463a <=( A167  and  A170 );
 a24467a <=( A200  and  A199 );
 a24468a <=( (not A166)  and  a24467a );
 a24469a <=( a24468a  and  a24463a );
 a24473a <=( A232  and  (not A202) );
 a24474a <=( (not A201)  and  a24473a );
 a24478a <=( A267  and  A266 );
 a24479a <=( A234  and  a24478a );
 a24480a <=( a24479a  and  a24474a );
 a24483a <=( A167  and  A170 );
 a24487a <=( A200  and  A199 );
 a24488a <=( (not A166)  and  a24487a );
 a24489a <=( a24488a  and  a24483a );
 a24493a <=( A233  and  (not A202) );
 a24494a <=( (not A201)  and  a24493a );
 a24498a <=( A300  and  A299 );
 a24499a <=( A234  and  a24498a );
 a24500a <=( a24499a  and  a24494a );
 a24503a <=( A167  and  A170 );
 a24507a <=( A200  and  A199 );
 a24508a <=( (not A166)  and  a24507a );
 a24509a <=( a24508a  and  a24503a );
 a24513a <=( A233  and  (not A202) );
 a24514a <=( (not A201)  and  a24513a );
 a24518a <=( A300  and  A298 );
 a24519a <=( A234  and  a24518a );
 a24520a <=( a24519a  and  a24514a );
 a24523a <=( A167  and  A170 );
 a24527a <=( A200  and  A199 );
 a24528a <=( (not A166)  and  a24527a );
 a24529a <=( a24528a  and  a24523a );
 a24533a <=( A233  and  (not A202) );
 a24534a <=( (not A201)  and  a24533a );
 a24538a <=( A267  and  A265 );
 a24539a <=( A234  and  a24538a );
 a24540a <=( a24539a  and  a24534a );
 a24543a <=( A167  and  A170 );
 a24547a <=( A200  and  A199 );
 a24548a <=( (not A166)  and  a24547a );
 a24549a <=( a24548a  and  a24543a );
 a24553a <=( A233  and  (not A202) );
 a24554a <=( (not A201)  and  a24553a );
 a24558a <=( A267  and  A266 );
 a24559a <=( A234  and  a24558a );
 a24560a <=( a24559a  and  a24554a );
 a24563a <=( A167  and  A170 );
 a24567a <=( A200  and  A199 );
 a24568a <=( (not A166)  and  a24567a );
 a24569a <=( a24568a  and  a24563a );
 a24573a <=( (not A232)  and  (not A202) );
 a24574a <=( (not A201)  and  a24573a );
 a24578a <=( A301  and  A236 );
 a24579a <=( A233  and  a24578a );
 a24580a <=( a24579a  and  a24574a );
 a24583a <=( A167  and  A170 );
 a24587a <=( A200  and  A199 );
 a24588a <=( (not A166)  and  a24587a );
 a24589a <=( a24588a  and  a24583a );
 a24593a <=( (not A232)  and  (not A202) );
 a24594a <=( (not A201)  and  a24593a );
 a24598a <=( A268  and  A236 );
 a24599a <=( A233  and  a24598a );
 a24600a <=( a24599a  and  a24594a );
 a24603a <=( A167  and  A170 );
 a24607a <=( A200  and  A199 );
 a24608a <=( (not A166)  and  a24607a );
 a24609a <=( a24608a  and  a24603a );
 a24613a <=( A232  and  (not A202) );
 a24614a <=( (not A201)  and  a24613a );
 a24618a <=( A301  and  A236 );
 a24619a <=( (not A233)  and  a24618a );
 a24620a <=( a24619a  and  a24614a );
 a24623a <=( A167  and  A170 );
 a24627a <=( A200  and  A199 );
 a24628a <=( (not A166)  and  a24627a );
 a24629a <=( a24628a  and  a24623a );
 a24633a <=( A232  and  (not A202) );
 a24634a <=( (not A201)  and  a24633a );
 a24638a <=( A268  and  A236 );
 a24639a <=( (not A233)  and  a24638a );
 a24640a <=( a24639a  and  a24634a );
 a24643a <=( A167  and  A170 );
 a24647a <=( (not A200)  and  (not A199) );
 a24648a <=( (not A166)  and  a24647a );
 a24649a <=( a24648a  and  a24643a );
 a24653a <=( A234  and  A232 );
 a24654a <=( (not A202)  and  a24653a );
 a24658a <=( A302  and  (not A299) );
 a24659a <=( A298  and  a24658a );
 a24660a <=( a24659a  and  a24654a );
 a24663a <=( A167  and  A170 );
 a24667a <=( (not A200)  and  (not A199) );
 a24668a <=( (not A166)  and  a24667a );
 a24669a <=( a24668a  and  a24663a );
 a24673a <=( A234  and  A232 );
 a24674a <=( (not A202)  and  a24673a );
 a24678a <=( A302  and  A299 );
 a24679a <=( (not A298)  and  a24678a );
 a24680a <=( a24679a  and  a24674a );
 a24683a <=( A167  and  A170 );
 a24687a <=( (not A200)  and  (not A199) );
 a24688a <=( (not A166)  and  a24687a );
 a24689a <=( a24688a  and  a24683a );
 a24693a <=( A234  and  A232 );
 a24694a <=( (not A202)  and  a24693a );
 a24698a <=( A269  and  A266 );
 a24699a <=( (not A265)  and  a24698a );
 a24700a <=( a24699a  and  a24694a );
 a24703a <=( A167  and  A170 );
 a24707a <=( (not A200)  and  (not A199) );
 a24708a <=( (not A166)  and  a24707a );
 a24709a <=( a24708a  and  a24703a );
 a24713a <=( A234  and  A232 );
 a24714a <=( (not A202)  and  a24713a );
 a24718a <=( A269  and  (not A266) );
 a24719a <=( A265  and  a24718a );
 a24720a <=( a24719a  and  a24714a );
 a24723a <=( A167  and  A170 );
 a24727a <=( (not A200)  and  (not A199) );
 a24728a <=( (not A166)  and  a24727a );
 a24729a <=( a24728a  and  a24723a );
 a24733a <=( A234  and  A233 );
 a24734a <=( (not A202)  and  a24733a );
 a24738a <=( A302  and  (not A299) );
 a24739a <=( A298  and  a24738a );
 a24740a <=( a24739a  and  a24734a );
 a24743a <=( A167  and  A170 );
 a24747a <=( (not A200)  and  (not A199) );
 a24748a <=( (not A166)  and  a24747a );
 a24749a <=( a24748a  and  a24743a );
 a24753a <=( A234  and  A233 );
 a24754a <=( (not A202)  and  a24753a );
 a24758a <=( A302  and  A299 );
 a24759a <=( (not A298)  and  a24758a );
 a24760a <=( a24759a  and  a24754a );
 a24763a <=( A167  and  A170 );
 a24767a <=( (not A200)  and  (not A199) );
 a24768a <=( (not A166)  and  a24767a );
 a24769a <=( a24768a  and  a24763a );
 a24773a <=( A234  and  A233 );
 a24774a <=( (not A202)  and  a24773a );
 a24778a <=( A269  and  A266 );
 a24779a <=( (not A265)  and  a24778a );
 a24780a <=( a24779a  and  a24774a );
 a24783a <=( A167  and  A170 );
 a24787a <=( (not A200)  and  (not A199) );
 a24788a <=( (not A166)  and  a24787a );
 a24789a <=( a24788a  and  a24783a );
 a24793a <=( A234  and  A233 );
 a24794a <=( (not A202)  and  a24793a );
 a24798a <=( A269  and  (not A266) );
 a24799a <=( A265  and  a24798a );
 a24800a <=( a24799a  and  a24794a );
 a24803a <=( A167  and  A170 );
 a24807a <=( (not A200)  and  (not A199) );
 a24808a <=( (not A166)  and  a24807a );
 a24809a <=( a24808a  and  a24803a );
 a24813a <=( A233  and  (not A232) );
 a24814a <=( (not A202)  and  a24813a );
 a24818a <=( A300  and  A299 );
 a24819a <=( A236  and  a24818a );
 a24820a <=( a24819a  and  a24814a );
 a24823a <=( A167  and  A170 );
 a24827a <=( (not A200)  and  (not A199) );
 a24828a <=( (not A166)  and  a24827a );
 a24829a <=( a24828a  and  a24823a );
 a24833a <=( A233  and  (not A232) );
 a24834a <=( (not A202)  and  a24833a );
 a24838a <=( A300  and  A298 );
 a24839a <=( A236  and  a24838a );
 a24840a <=( a24839a  and  a24834a );
 a24843a <=( A167  and  A170 );
 a24847a <=( (not A200)  and  (not A199) );
 a24848a <=( (not A166)  and  a24847a );
 a24849a <=( a24848a  and  a24843a );
 a24853a <=( A233  and  (not A232) );
 a24854a <=( (not A202)  and  a24853a );
 a24858a <=( A267  and  A265 );
 a24859a <=( A236  and  a24858a );
 a24860a <=( a24859a  and  a24854a );
 a24863a <=( A167  and  A170 );
 a24867a <=( (not A200)  and  (not A199) );
 a24868a <=( (not A166)  and  a24867a );
 a24869a <=( a24868a  and  a24863a );
 a24873a <=( A233  and  (not A232) );
 a24874a <=( (not A202)  and  a24873a );
 a24878a <=( A267  and  A266 );
 a24879a <=( A236  and  a24878a );
 a24880a <=( a24879a  and  a24874a );
 a24883a <=( A167  and  A170 );
 a24887a <=( (not A200)  and  (not A199) );
 a24888a <=( (not A166)  and  a24887a );
 a24889a <=( a24888a  and  a24883a );
 a24893a <=( (not A233)  and  A232 );
 a24894a <=( (not A202)  and  a24893a );
 a24898a <=( A300  and  A299 );
 a24899a <=( A236  and  a24898a );
 a24900a <=( a24899a  and  a24894a );
 a24903a <=( A167  and  A170 );
 a24907a <=( (not A200)  and  (not A199) );
 a24908a <=( (not A166)  and  a24907a );
 a24909a <=( a24908a  and  a24903a );
 a24913a <=( (not A233)  and  A232 );
 a24914a <=( (not A202)  and  a24913a );
 a24918a <=( A300  and  A298 );
 a24919a <=( A236  and  a24918a );
 a24920a <=( a24919a  and  a24914a );
 a24923a <=( A167  and  A170 );
 a24927a <=( (not A200)  and  (not A199) );
 a24928a <=( (not A166)  and  a24927a );
 a24929a <=( a24928a  and  a24923a );
 a24933a <=( (not A233)  and  A232 );
 a24934a <=( (not A202)  and  a24933a );
 a24938a <=( A267  and  A265 );
 a24939a <=( A236  and  a24938a );
 a24940a <=( a24939a  and  a24934a );
 a24943a <=( A167  and  A170 );
 a24947a <=( (not A200)  and  (not A199) );
 a24948a <=( (not A166)  and  a24947a );
 a24949a <=( a24948a  and  a24943a );
 a24953a <=( (not A233)  and  A232 );
 a24954a <=( (not A202)  and  a24953a );
 a24958a <=( A267  and  A266 );
 a24959a <=( A236  and  a24958a );
 a24960a <=( a24959a  and  a24954a );
 a24963a <=( (not A167)  and  A170 );
 a24967a <=( (not A202)  and  (not A201) );
 a24968a <=( A166  and  a24967a );
 a24969a <=( a24968a  and  a24963a );
 a24973a <=( A234  and  A232 );
 a24974a <=( (not A203)  and  a24973a );
 a24978a <=( A302  and  (not A299) );
 a24979a <=( A298  and  a24978a );
 a24980a <=( a24979a  and  a24974a );
 a24983a <=( (not A167)  and  A170 );
 a24987a <=( (not A202)  and  (not A201) );
 a24988a <=( A166  and  a24987a );
 a24989a <=( a24988a  and  a24983a );
 a24993a <=( A234  and  A232 );
 a24994a <=( (not A203)  and  a24993a );
 a24998a <=( A302  and  A299 );
 a24999a <=( (not A298)  and  a24998a );
 a25000a <=( a24999a  and  a24994a );
 a25003a <=( (not A167)  and  A170 );
 a25007a <=( (not A202)  and  (not A201) );
 a25008a <=( A166  and  a25007a );
 a25009a <=( a25008a  and  a25003a );
 a25013a <=( A234  and  A232 );
 a25014a <=( (not A203)  and  a25013a );
 a25018a <=( A269  and  A266 );
 a25019a <=( (not A265)  and  a25018a );
 a25020a <=( a25019a  and  a25014a );
 a25023a <=( (not A167)  and  A170 );
 a25027a <=( (not A202)  and  (not A201) );
 a25028a <=( A166  and  a25027a );
 a25029a <=( a25028a  and  a25023a );
 a25033a <=( A234  and  A232 );
 a25034a <=( (not A203)  and  a25033a );
 a25038a <=( A269  and  (not A266) );
 a25039a <=( A265  and  a25038a );
 a25040a <=( a25039a  and  a25034a );
 a25043a <=( (not A167)  and  A170 );
 a25047a <=( (not A202)  and  (not A201) );
 a25048a <=( A166  and  a25047a );
 a25049a <=( a25048a  and  a25043a );
 a25053a <=( A234  and  A233 );
 a25054a <=( (not A203)  and  a25053a );
 a25058a <=( A302  and  (not A299) );
 a25059a <=( A298  and  a25058a );
 a25060a <=( a25059a  and  a25054a );
 a25063a <=( (not A167)  and  A170 );
 a25067a <=( (not A202)  and  (not A201) );
 a25068a <=( A166  and  a25067a );
 a25069a <=( a25068a  and  a25063a );
 a25073a <=( A234  and  A233 );
 a25074a <=( (not A203)  and  a25073a );
 a25078a <=( A302  and  A299 );
 a25079a <=( (not A298)  and  a25078a );
 a25080a <=( a25079a  and  a25074a );
 a25083a <=( (not A167)  and  A170 );
 a25087a <=( (not A202)  and  (not A201) );
 a25088a <=( A166  and  a25087a );
 a25089a <=( a25088a  and  a25083a );
 a25093a <=( A234  and  A233 );
 a25094a <=( (not A203)  and  a25093a );
 a25098a <=( A269  and  A266 );
 a25099a <=( (not A265)  and  a25098a );
 a25100a <=( a25099a  and  a25094a );
 a25103a <=( (not A167)  and  A170 );
 a25107a <=( (not A202)  and  (not A201) );
 a25108a <=( A166  and  a25107a );
 a25109a <=( a25108a  and  a25103a );
 a25113a <=( A234  and  A233 );
 a25114a <=( (not A203)  and  a25113a );
 a25118a <=( A269  and  (not A266) );
 a25119a <=( A265  and  a25118a );
 a25120a <=( a25119a  and  a25114a );
 a25123a <=( (not A167)  and  A170 );
 a25127a <=( (not A202)  and  (not A201) );
 a25128a <=( A166  and  a25127a );
 a25129a <=( a25128a  and  a25123a );
 a25133a <=( A233  and  (not A232) );
 a25134a <=( (not A203)  and  a25133a );
 a25138a <=( A300  and  A299 );
 a25139a <=( A236  and  a25138a );
 a25140a <=( a25139a  and  a25134a );
 a25143a <=( (not A167)  and  A170 );
 a25147a <=( (not A202)  and  (not A201) );
 a25148a <=( A166  and  a25147a );
 a25149a <=( a25148a  and  a25143a );
 a25153a <=( A233  and  (not A232) );
 a25154a <=( (not A203)  and  a25153a );
 a25158a <=( A300  and  A298 );
 a25159a <=( A236  and  a25158a );
 a25160a <=( a25159a  and  a25154a );
 a25163a <=( (not A167)  and  A170 );
 a25167a <=( (not A202)  and  (not A201) );
 a25168a <=( A166  and  a25167a );
 a25169a <=( a25168a  and  a25163a );
 a25173a <=( A233  and  (not A232) );
 a25174a <=( (not A203)  and  a25173a );
 a25178a <=( A267  and  A265 );
 a25179a <=( A236  and  a25178a );
 a25180a <=( a25179a  and  a25174a );
 a25183a <=( (not A167)  and  A170 );
 a25187a <=( (not A202)  and  (not A201) );
 a25188a <=( A166  and  a25187a );
 a25189a <=( a25188a  and  a25183a );
 a25193a <=( A233  and  (not A232) );
 a25194a <=( (not A203)  and  a25193a );
 a25198a <=( A267  and  A266 );
 a25199a <=( A236  and  a25198a );
 a25200a <=( a25199a  and  a25194a );
 a25203a <=( (not A167)  and  A170 );
 a25207a <=( (not A202)  and  (not A201) );
 a25208a <=( A166  and  a25207a );
 a25209a <=( a25208a  and  a25203a );
 a25213a <=( (not A233)  and  A232 );
 a25214a <=( (not A203)  and  a25213a );
 a25218a <=( A300  and  A299 );
 a25219a <=( A236  and  a25218a );
 a25220a <=( a25219a  and  a25214a );
 a25223a <=( (not A167)  and  A170 );
 a25227a <=( (not A202)  and  (not A201) );
 a25228a <=( A166  and  a25227a );
 a25229a <=( a25228a  and  a25223a );
 a25233a <=( (not A233)  and  A232 );
 a25234a <=( (not A203)  and  a25233a );
 a25238a <=( A300  and  A298 );
 a25239a <=( A236  and  a25238a );
 a25240a <=( a25239a  and  a25234a );
 a25243a <=( (not A167)  and  A170 );
 a25247a <=( (not A202)  and  (not A201) );
 a25248a <=( A166  and  a25247a );
 a25249a <=( a25248a  and  a25243a );
 a25253a <=( (not A233)  and  A232 );
 a25254a <=( (not A203)  and  a25253a );
 a25258a <=( A267  and  A265 );
 a25259a <=( A236  and  a25258a );
 a25260a <=( a25259a  and  a25254a );
 a25263a <=( (not A167)  and  A170 );
 a25267a <=( (not A202)  and  (not A201) );
 a25268a <=( A166  and  a25267a );
 a25269a <=( a25268a  and  a25263a );
 a25273a <=( (not A233)  and  A232 );
 a25274a <=( (not A203)  and  a25273a );
 a25278a <=( A267  and  A266 );
 a25279a <=( A236  and  a25278a );
 a25280a <=( a25279a  and  a25274a );
 a25283a <=( (not A167)  and  A170 );
 a25287a <=( A200  and  A199 );
 a25288a <=( A166  and  a25287a );
 a25289a <=( a25288a  and  a25283a );
 a25293a <=( A235  and  (not A202) );
 a25294a <=( (not A201)  and  a25293a );
 a25298a <=( A302  and  (not A299) );
 a25299a <=( A298  and  a25298a );
 a25300a <=( a25299a  and  a25294a );
 a25303a <=( (not A167)  and  A170 );
 a25307a <=( A200  and  A199 );
 a25308a <=( A166  and  a25307a );
 a25309a <=( a25308a  and  a25303a );
 a25313a <=( A235  and  (not A202) );
 a25314a <=( (not A201)  and  a25313a );
 a25318a <=( A302  and  A299 );
 a25319a <=( (not A298)  and  a25318a );
 a25320a <=( a25319a  and  a25314a );
 a25323a <=( (not A167)  and  A170 );
 a25327a <=( A200  and  A199 );
 a25328a <=( A166  and  a25327a );
 a25329a <=( a25328a  and  a25323a );
 a25333a <=( A235  and  (not A202) );
 a25334a <=( (not A201)  and  a25333a );
 a25338a <=( A269  and  A266 );
 a25339a <=( (not A265)  and  a25338a );
 a25340a <=( a25339a  and  a25334a );
 a25343a <=( (not A167)  and  A170 );
 a25347a <=( A200  and  A199 );
 a25348a <=( A166  and  a25347a );
 a25349a <=( a25348a  and  a25343a );
 a25353a <=( A235  and  (not A202) );
 a25354a <=( (not A201)  and  a25353a );
 a25358a <=( A269  and  (not A266) );
 a25359a <=( A265  and  a25358a );
 a25360a <=( a25359a  and  a25354a );
 a25363a <=( (not A167)  and  A170 );
 a25367a <=( A200  and  A199 );
 a25368a <=( A166  and  a25367a );
 a25369a <=( a25368a  and  a25363a );
 a25373a <=( A232  and  (not A202) );
 a25374a <=( (not A201)  and  a25373a );
 a25378a <=( A300  and  A299 );
 a25379a <=( A234  and  a25378a );
 a25380a <=( a25379a  and  a25374a );
 a25383a <=( (not A167)  and  A170 );
 a25387a <=( A200  and  A199 );
 a25388a <=( A166  and  a25387a );
 a25389a <=( a25388a  and  a25383a );
 a25393a <=( A232  and  (not A202) );
 a25394a <=( (not A201)  and  a25393a );
 a25398a <=( A300  and  A298 );
 a25399a <=( A234  and  a25398a );
 a25400a <=( a25399a  and  a25394a );
 a25403a <=( (not A167)  and  A170 );
 a25407a <=( A200  and  A199 );
 a25408a <=( A166  and  a25407a );
 a25409a <=( a25408a  and  a25403a );
 a25413a <=( A232  and  (not A202) );
 a25414a <=( (not A201)  and  a25413a );
 a25418a <=( A267  and  A265 );
 a25419a <=( A234  and  a25418a );
 a25420a <=( a25419a  and  a25414a );
 a25423a <=( (not A167)  and  A170 );
 a25427a <=( A200  and  A199 );
 a25428a <=( A166  and  a25427a );
 a25429a <=( a25428a  and  a25423a );
 a25433a <=( A232  and  (not A202) );
 a25434a <=( (not A201)  and  a25433a );
 a25438a <=( A267  and  A266 );
 a25439a <=( A234  and  a25438a );
 a25440a <=( a25439a  and  a25434a );
 a25443a <=( (not A167)  and  A170 );
 a25447a <=( A200  and  A199 );
 a25448a <=( A166  and  a25447a );
 a25449a <=( a25448a  and  a25443a );
 a25453a <=( A233  and  (not A202) );
 a25454a <=( (not A201)  and  a25453a );
 a25458a <=( A300  and  A299 );
 a25459a <=( A234  and  a25458a );
 a25460a <=( a25459a  and  a25454a );
 a25463a <=( (not A167)  and  A170 );
 a25467a <=( A200  and  A199 );
 a25468a <=( A166  and  a25467a );
 a25469a <=( a25468a  and  a25463a );
 a25473a <=( A233  and  (not A202) );
 a25474a <=( (not A201)  and  a25473a );
 a25478a <=( A300  and  A298 );
 a25479a <=( A234  and  a25478a );
 a25480a <=( a25479a  and  a25474a );
 a25483a <=( (not A167)  and  A170 );
 a25487a <=( A200  and  A199 );
 a25488a <=( A166  and  a25487a );
 a25489a <=( a25488a  and  a25483a );
 a25493a <=( A233  and  (not A202) );
 a25494a <=( (not A201)  and  a25493a );
 a25498a <=( A267  and  A265 );
 a25499a <=( A234  and  a25498a );
 a25500a <=( a25499a  and  a25494a );
 a25503a <=( (not A167)  and  A170 );
 a25507a <=( A200  and  A199 );
 a25508a <=( A166  and  a25507a );
 a25509a <=( a25508a  and  a25503a );
 a25513a <=( A233  and  (not A202) );
 a25514a <=( (not A201)  and  a25513a );
 a25518a <=( A267  and  A266 );
 a25519a <=( A234  and  a25518a );
 a25520a <=( a25519a  and  a25514a );
 a25523a <=( (not A167)  and  A170 );
 a25527a <=( A200  and  A199 );
 a25528a <=( A166  and  a25527a );
 a25529a <=( a25528a  and  a25523a );
 a25533a <=( (not A232)  and  (not A202) );
 a25534a <=( (not A201)  and  a25533a );
 a25538a <=( A301  and  A236 );
 a25539a <=( A233  and  a25538a );
 a25540a <=( a25539a  and  a25534a );
 a25543a <=( (not A167)  and  A170 );
 a25547a <=( A200  and  A199 );
 a25548a <=( A166  and  a25547a );
 a25549a <=( a25548a  and  a25543a );
 a25553a <=( (not A232)  and  (not A202) );
 a25554a <=( (not A201)  and  a25553a );
 a25558a <=( A268  and  A236 );
 a25559a <=( A233  and  a25558a );
 a25560a <=( a25559a  and  a25554a );
 a25563a <=( (not A167)  and  A170 );
 a25567a <=( A200  and  A199 );
 a25568a <=( A166  and  a25567a );
 a25569a <=( a25568a  and  a25563a );
 a25573a <=( A232  and  (not A202) );
 a25574a <=( (not A201)  and  a25573a );
 a25578a <=( A301  and  A236 );
 a25579a <=( (not A233)  and  a25578a );
 a25580a <=( a25579a  and  a25574a );
 a25583a <=( (not A167)  and  A170 );
 a25587a <=( A200  and  A199 );
 a25588a <=( A166  and  a25587a );
 a25589a <=( a25588a  and  a25583a );
 a25593a <=( A232  and  (not A202) );
 a25594a <=( (not A201)  and  a25593a );
 a25598a <=( A268  and  A236 );
 a25599a <=( (not A233)  and  a25598a );
 a25600a <=( a25599a  and  a25594a );
 a25603a <=( (not A167)  and  A170 );
 a25607a <=( (not A200)  and  (not A199) );
 a25608a <=( A166  and  a25607a );
 a25609a <=( a25608a  and  a25603a );
 a25613a <=( A234  and  A232 );
 a25614a <=( (not A202)  and  a25613a );
 a25618a <=( A302  and  (not A299) );
 a25619a <=( A298  and  a25618a );
 a25620a <=( a25619a  and  a25614a );
 a25623a <=( (not A167)  and  A170 );
 a25627a <=( (not A200)  and  (not A199) );
 a25628a <=( A166  and  a25627a );
 a25629a <=( a25628a  and  a25623a );
 a25633a <=( A234  and  A232 );
 a25634a <=( (not A202)  and  a25633a );
 a25638a <=( A302  and  A299 );
 a25639a <=( (not A298)  and  a25638a );
 a25640a <=( a25639a  and  a25634a );
 a25643a <=( (not A167)  and  A170 );
 a25647a <=( (not A200)  and  (not A199) );
 a25648a <=( A166  and  a25647a );
 a25649a <=( a25648a  and  a25643a );
 a25653a <=( A234  and  A232 );
 a25654a <=( (not A202)  and  a25653a );
 a25658a <=( A269  and  A266 );
 a25659a <=( (not A265)  and  a25658a );
 a25660a <=( a25659a  and  a25654a );
 a25663a <=( (not A167)  and  A170 );
 a25667a <=( (not A200)  and  (not A199) );
 a25668a <=( A166  and  a25667a );
 a25669a <=( a25668a  and  a25663a );
 a25673a <=( A234  and  A232 );
 a25674a <=( (not A202)  and  a25673a );
 a25678a <=( A269  and  (not A266) );
 a25679a <=( A265  and  a25678a );
 a25680a <=( a25679a  and  a25674a );
 a25683a <=( (not A167)  and  A170 );
 a25687a <=( (not A200)  and  (not A199) );
 a25688a <=( A166  and  a25687a );
 a25689a <=( a25688a  and  a25683a );
 a25693a <=( A234  and  A233 );
 a25694a <=( (not A202)  and  a25693a );
 a25698a <=( A302  and  (not A299) );
 a25699a <=( A298  and  a25698a );
 a25700a <=( a25699a  and  a25694a );
 a25703a <=( (not A167)  and  A170 );
 a25707a <=( (not A200)  and  (not A199) );
 a25708a <=( A166  and  a25707a );
 a25709a <=( a25708a  and  a25703a );
 a25713a <=( A234  and  A233 );
 a25714a <=( (not A202)  and  a25713a );
 a25718a <=( A302  and  A299 );
 a25719a <=( (not A298)  and  a25718a );
 a25720a <=( a25719a  and  a25714a );
 a25723a <=( (not A167)  and  A170 );
 a25727a <=( (not A200)  and  (not A199) );
 a25728a <=( A166  and  a25727a );
 a25729a <=( a25728a  and  a25723a );
 a25733a <=( A234  and  A233 );
 a25734a <=( (not A202)  and  a25733a );
 a25738a <=( A269  and  A266 );
 a25739a <=( (not A265)  and  a25738a );
 a25740a <=( a25739a  and  a25734a );
 a25743a <=( (not A167)  and  A170 );
 a25747a <=( (not A200)  and  (not A199) );
 a25748a <=( A166  and  a25747a );
 a25749a <=( a25748a  and  a25743a );
 a25753a <=( A234  and  A233 );
 a25754a <=( (not A202)  and  a25753a );
 a25758a <=( A269  and  (not A266) );
 a25759a <=( A265  and  a25758a );
 a25760a <=( a25759a  and  a25754a );
 a25763a <=( (not A167)  and  A170 );
 a25767a <=( (not A200)  and  (not A199) );
 a25768a <=( A166  and  a25767a );
 a25769a <=( a25768a  and  a25763a );
 a25773a <=( A233  and  (not A232) );
 a25774a <=( (not A202)  and  a25773a );
 a25778a <=( A300  and  A299 );
 a25779a <=( A236  and  a25778a );
 a25780a <=( a25779a  and  a25774a );
 a25783a <=( (not A167)  and  A170 );
 a25787a <=( (not A200)  and  (not A199) );
 a25788a <=( A166  and  a25787a );
 a25789a <=( a25788a  and  a25783a );
 a25793a <=( A233  and  (not A232) );
 a25794a <=( (not A202)  and  a25793a );
 a25798a <=( A300  and  A298 );
 a25799a <=( A236  and  a25798a );
 a25800a <=( a25799a  and  a25794a );
 a25803a <=( (not A167)  and  A170 );
 a25807a <=( (not A200)  and  (not A199) );
 a25808a <=( A166  and  a25807a );
 a25809a <=( a25808a  and  a25803a );
 a25813a <=( A233  and  (not A232) );
 a25814a <=( (not A202)  and  a25813a );
 a25818a <=( A267  and  A265 );
 a25819a <=( A236  and  a25818a );
 a25820a <=( a25819a  and  a25814a );
 a25823a <=( (not A167)  and  A170 );
 a25827a <=( (not A200)  and  (not A199) );
 a25828a <=( A166  and  a25827a );
 a25829a <=( a25828a  and  a25823a );
 a25833a <=( A233  and  (not A232) );
 a25834a <=( (not A202)  and  a25833a );
 a25838a <=( A267  and  A266 );
 a25839a <=( A236  and  a25838a );
 a25840a <=( a25839a  and  a25834a );
 a25843a <=( (not A167)  and  A170 );
 a25847a <=( (not A200)  and  (not A199) );
 a25848a <=( A166  and  a25847a );
 a25849a <=( a25848a  and  a25843a );
 a25853a <=( (not A233)  and  A232 );
 a25854a <=( (not A202)  and  a25853a );
 a25858a <=( A300  and  A299 );
 a25859a <=( A236  and  a25858a );
 a25860a <=( a25859a  and  a25854a );
 a25863a <=( (not A167)  and  A170 );
 a25867a <=( (not A200)  and  (not A199) );
 a25868a <=( A166  and  a25867a );
 a25869a <=( a25868a  and  a25863a );
 a25873a <=( (not A233)  and  A232 );
 a25874a <=( (not A202)  and  a25873a );
 a25878a <=( A300  and  A298 );
 a25879a <=( A236  and  a25878a );
 a25880a <=( a25879a  and  a25874a );
 a25883a <=( (not A167)  and  A170 );
 a25887a <=( (not A200)  and  (not A199) );
 a25888a <=( A166  and  a25887a );
 a25889a <=( a25888a  and  a25883a );
 a25893a <=( (not A233)  and  A232 );
 a25894a <=( (not A202)  and  a25893a );
 a25898a <=( A267  and  A265 );
 a25899a <=( A236  and  a25898a );
 a25900a <=( a25899a  and  a25894a );
 a25903a <=( (not A167)  and  A170 );
 a25907a <=( (not A200)  and  (not A199) );
 a25908a <=( A166  and  a25907a );
 a25909a <=( a25908a  and  a25903a );
 a25913a <=( (not A233)  and  A232 );
 a25914a <=( (not A202)  and  a25913a );
 a25918a <=( A267  and  A266 );
 a25919a <=( A236  and  a25918a );
 a25920a <=( a25919a  and  a25914a );
 a25923a <=( A199  and  A169 );
 a25927a <=( (not A202)  and  (not A201) );
 a25928a <=( A200  and  a25927a );
 a25929a <=( a25928a  and  a25923a );
 a25933a <=( A236  and  A233 );
 a25934a <=( (not A232)  and  a25933a );
 a25938a <=( A302  and  (not A299) );
 a25939a <=( A298  and  a25938a );
 a25940a <=( a25939a  and  a25934a );
 a25943a <=( A199  and  A169 );
 a25947a <=( (not A202)  and  (not A201) );
 a25948a <=( A200  and  a25947a );
 a25949a <=( a25948a  and  a25943a );
 a25953a <=( A236  and  A233 );
 a25954a <=( (not A232)  and  a25953a );
 a25958a <=( A302  and  A299 );
 a25959a <=( (not A298)  and  a25958a );
 a25960a <=( a25959a  and  a25954a );
 a25963a <=( A199  and  A169 );
 a25967a <=( (not A202)  and  (not A201) );
 a25968a <=( A200  and  a25967a );
 a25969a <=( a25968a  and  a25963a );
 a25973a <=( A236  and  A233 );
 a25974a <=( (not A232)  and  a25973a );
 a25978a <=( A269  and  A266 );
 a25979a <=( (not A265)  and  a25978a );
 a25980a <=( a25979a  and  a25974a );
 a25983a <=( A199  and  A169 );
 a25987a <=( (not A202)  and  (not A201) );
 a25988a <=( A200  and  a25987a );
 a25989a <=( a25988a  and  a25983a );
 a25993a <=( A236  and  A233 );
 a25994a <=( (not A232)  and  a25993a );
 a25998a <=( A269  and  (not A266) );
 a25999a <=( A265  and  a25998a );
 a26000a <=( a25999a  and  a25994a );
 a26003a <=( A199  and  A169 );
 a26007a <=( (not A202)  and  (not A201) );
 a26008a <=( A200  and  a26007a );
 a26009a <=( a26008a  and  a26003a );
 a26013a <=( A236  and  (not A233) );
 a26014a <=( A232  and  a26013a );
 a26018a <=( A302  and  (not A299) );
 a26019a <=( A298  and  a26018a );
 a26020a <=( a26019a  and  a26014a );
 a26023a <=( A199  and  A169 );
 a26027a <=( (not A202)  and  (not A201) );
 a26028a <=( A200  and  a26027a );
 a26029a <=( a26028a  and  a26023a );
 a26033a <=( A236  and  (not A233) );
 a26034a <=( A232  and  a26033a );
 a26038a <=( A302  and  A299 );
 a26039a <=( (not A298)  and  a26038a );
 a26040a <=( a26039a  and  a26034a );
 a26043a <=( A199  and  A169 );
 a26047a <=( (not A202)  and  (not A201) );
 a26048a <=( A200  and  a26047a );
 a26049a <=( a26048a  and  a26043a );
 a26053a <=( A236  and  (not A233) );
 a26054a <=( A232  and  a26053a );
 a26058a <=( A269  and  A266 );
 a26059a <=( (not A265)  and  a26058a );
 a26060a <=( a26059a  and  a26054a );
 a26063a <=( A199  and  A169 );
 a26067a <=( (not A202)  and  (not A201) );
 a26068a <=( A200  and  a26067a );
 a26069a <=( a26068a  and  a26063a );
 a26073a <=( A236  and  (not A233) );
 a26074a <=( A232  and  a26073a );
 a26078a <=( A269  and  (not A266) );
 a26079a <=( A265  and  a26078a );
 a26080a <=( a26079a  and  a26074a );
 a26083a <=( (not A167)  and  (not A169) );
 a26087a <=( A201  and  A199 );
 a26088a <=( (not A166)  and  a26087a );
 a26089a <=( a26088a  and  a26083a );
 a26093a <=( A236  and  A233 );
 a26094a <=( (not A232)  and  a26093a );
 a26098a <=( A302  and  (not A299) );
 a26099a <=( A298  and  a26098a );
 a26100a <=( a26099a  and  a26094a );
 a26103a <=( (not A167)  and  (not A169) );
 a26107a <=( A201  and  A199 );
 a26108a <=( (not A166)  and  a26107a );
 a26109a <=( a26108a  and  a26103a );
 a26113a <=( A236  and  A233 );
 a26114a <=( (not A232)  and  a26113a );
 a26118a <=( A302  and  A299 );
 a26119a <=( (not A298)  and  a26118a );
 a26120a <=( a26119a  and  a26114a );
 a26123a <=( (not A167)  and  (not A169) );
 a26127a <=( A201  and  A199 );
 a26128a <=( (not A166)  and  a26127a );
 a26129a <=( a26128a  and  a26123a );
 a26133a <=( A236  and  A233 );
 a26134a <=( (not A232)  and  a26133a );
 a26138a <=( A269  and  A266 );
 a26139a <=( (not A265)  and  a26138a );
 a26140a <=( a26139a  and  a26134a );
 a26143a <=( (not A167)  and  (not A169) );
 a26147a <=( A201  and  A199 );
 a26148a <=( (not A166)  and  a26147a );
 a26149a <=( a26148a  and  a26143a );
 a26153a <=( A236  and  A233 );
 a26154a <=( (not A232)  and  a26153a );
 a26158a <=( A269  and  (not A266) );
 a26159a <=( A265  and  a26158a );
 a26160a <=( a26159a  and  a26154a );
 a26163a <=( (not A167)  and  (not A169) );
 a26167a <=( A201  and  A199 );
 a26168a <=( (not A166)  and  a26167a );
 a26169a <=( a26168a  and  a26163a );
 a26173a <=( A236  and  (not A233) );
 a26174a <=( A232  and  a26173a );
 a26178a <=( A302  and  (not A299) );
 a26179a <=( A298  and  a26178a );
 a26180a <=( a26179a  and  a26174a );
 a26183a <=( (not A167)  and  (not A169) );
 a26187a <=( A201  and  A199 );
 a26188a <=( (not A166)  and  a26187a );
 a26189a <=( a26188a  and  a26183a );
 a26193a <=( A236  and  (not A233) );
 a26194a <=( A232  and  a26193a );
 a26198a <=( A302  and  A299 );
 a26199a <=( (not A298)  and  a26198a );
 a26200a <=( a26199a  and  a26194a );
 a26203a <=( (not A167)  and  (not A169) );
 a26207a <=( A201  and  A199 );
 a26208a <=( (not A166)  and  a26207a );
 a26209a <=( a26208a  and  a26203a );
 a26213a <=( A236  and  (not A233) );
 a26214a <=( A232  and  a26213a );
 a26218a <=( A269  and  A266 );
 a26219a <=( (not A265)  and  a26218a );
 a26220a <=( a26219a  and  a26214a );
 a26223a <=( (not A167)  and  (not A169) );
 a26227a <=( A201  and  A199 );
 a26228a <=( (not A166)  and  a26227a );
 a26229a <=( a26228a  and  a26223a );
 a26233a <=( A236  and  (not A233) );
 a26234a <=( A232  and  a26233a );
 a26238a <=( A269  and  (not A266) );
 a26239a <=( A265  and  a26238a );
 a26240a <=( a26239a  and  a26234a );
 a26243a <=( (not A167)  and  (not A169) );
 a26247a <=( A201  and  A200 );
 a26248a <=( (not A166)  and  a26247a );
 a26249a <=( a26248a  and  a26243a );
 a26253a <=( A236  and  A233 );
 a26254a <=( (not A232)  and  a26253a );
 a26258a <=( A302  and  (not A299) );
 a26259a <=( A298  and  a26258a );
 a26260a <=( a26259a  and  a26254a );
 a26263a <=( (not A167)  and  (not A169) );
 a26267a <=( A201  and  A200 );
 a26268a <=( (not A166)  and  a26267a );
 a26269a <=( a26268a  and  a26263a );
 a26273a <=( A236  and  A233 );
 a26274a <=( (not A232)  and  a26273a );
 a26278a <=( A302  and  A299 );
 a26279a <=( (not A298)  and  a26278a );
 a26280a <=( a26279a  and  a26274a );
 a26283a <=( (not A167)  and  (not A169) );
 a26287a <=( A201  and  A200 );
 a26288a <=( (not A166)  and  a26287a );
 a26289a <=( a26288a  and  a26283a );
 a26293a <=( A236  and  A233 );
 a26294a <=( (not A232)  and  a26293a );
 a26298a <=( A269  and  A266 );
 a26299a <=( (not A265)  and  a26298a );
 a26300a <=( a26299a  and  a26294a );
 a26303a <=( (not A167)  and  (not A169) );
 a26307a <=( A201  and  A200 );
 a26308a <=( (not A166)  and  a26307a );
 a26309a <=( a26308a  and  a26303a );
 a26313a <=( A236  and  A233 );
 a26314a <=( (not A232)  and  a26313a );
 a26318a <=( A269  and  (not A266) );
 a26319a <=( A265  and  a26318a );
 a26320a <=( a26319a  and  a26314a );
 a26323a <=( (not A167)  and  (not A169) );
 a26327a <=( A201  and  A200 );
 a26328a <=( (not A166)  and  a26327a );
 a26329a <=( a26328a  and  a26323a );
 a26333a <=( A236  and  (not A233) );
 a26334a <=( A232  and  a26333a );
 a26338a <=( A302  and  (not A299) );
 a26339a <=( A298  and  a26338a );
 a26340a <=( a26339a  and  a26334a );
 a26343a <=( (not A167)  and  (not A169) );
 a26347a <=( A201  and  A200 );
 a26348a <=( (not A166)  and  a26347a );
 a26349a <=( a26348a  and  a26343a );
 a26353a <=( A236  and  (not A233) );
 a26354a <=( A232  and  a26353a );
 a26358a <=( A302  and  A299 );
 a26359a <=( (not A298)  and  a26358a );
 a26360a <=( a26359a  and  a26354a );
 a26363a <=( (not A167)  and  (not A169) );
 a26367a <=( A201  and  A200 );
 a26368a <=( (not A166)  and  a26367a );
 a26369a <=( a26368a  and  a26363a );
 a26373a <=( A236  and  (not A233) );
 a26374a <=( A232  and  a26373a );
 a26378a <=( A269  and  A266 );
 a26379a <=( (not A265)  and  a26378a );
 a26380a <=( a26379a  and  a26374a );
 a26383a <=( (not A167)  and  (not A169) );
 a26387a <=( A201  and  A200 );
 a26388a <=( (not A166)  and  a26387a );
 a26389a <=( a26388a  and  a26383a );
 a26393a <=( A236  and  (not A233) );
 a26394a <=( A232  and  a26393a );
 a26398a <=( A269  and  (not A266) );
 a26399a <=( A265  and  a26398a );
 a26400a <=( a26399a  and  a26394a );
 a26403a <=( (not A167)  and  (not A169) );
 a26407a <=( A200  and  (not A199) );
 a26408a <=( (not A166)  and  a26407a );
 a26409a <=( a26408a  and  a26403a );
 a26413a <=( A234  and  A232 );
 a26414a <=( A203  and  a26413a );
 a26418a <=( A302  and  (not A299) );
 a26419a <=( A298  and  a26418a );
 a26420a <=( a26419a  and  a26414a );
 a26423a <=( (not A167)  and  (not A169) );
 a26427a <=( A200  and  (not A199) );
 a26428a <=( (not A166)  and  a26427a );
 a26429a <=( a26428a  and  a26423a );
 a26433a <=( A234  and  A232 );
 a26434a <=( A203  and  a26433a );
 a26438a <=( A302  and  A299 );
 a26439a <=( (not A298)  and  a26438a );
 a26440a <=( a26439a  and  a26434a );
 a26443a <=( (not A167)  and  (not A169) );
 a26447a <=( A200  and  (not A199) );
 a26448a <=( (not A166)  and  a26447a );
 a26449a <=( a26448a  and  a26443a );
 a26453a <=( A234  and  A232 );
 a26454a <=( A203  and  a26453a );
 a26458a <=( A269  and  A266 );
 a26459a <=( (not A265)  and  a26458a );
 a26460a <=( a26459a  and  a26454a );
 a26463a <=( (not A167)  and  (not A169) );
 a26467a <=( A200  and  (not A199) );
 a26468a <=( (not A166)  and  a26467a );
 a26469a <=( a26468a  and  a26463a );
 a26473a <=( A234  and  A232 );
 a26474a <=( A203  and  a26473a );
 a26478a <=( A269  and  (not A266) );
 a26479a <=( A265  and  a26478a );
 a26480a <=( a26479a  and  a26474a );
 a26483a <=( (not A167)  and  (not A169) );
 a26487a <=( A200  and  (not A199) );
 a26488a <=( (not A166)  and  a26487a );
 a26489a <=( a26488a  and  a26483a );
 a26493a <=( A234  and  A233 );
 a26494a <=( A203  and  a26493a );
 a26498a <=( A302  and  (not A299) );
 a26499a <=( A298  and  a26498a );
 a26500a <=( a26499a  and  a26494a );
 a26503a <=( (not A167)  and  (not A169) );
 a26507a <=( A200  and  (not A199) );
 a26508a <=( (not A166)  and  a26507a );
 a26509a <=( a26508a  and  a26503a );
 a26513a <=( A234  and  A233 );
 a26514a <=( A203  and  a26513a );
 a26518a <=( A302  and  A299 );
 a26519a <=( (not A298)  and  a26518a );
 a26520a <=( a26519a  and  a26514a );
 a26523a <=( (not A167)  and  (not A169) );
 a26527a <=( A200  and  (not A199) );
 a26528a <=( (not A166)  and  a26527a );
 a26529a <=( a26528a  and  a26523a );
 a26533a <=( A234  and  A233 );
 a26534a <=( A203  and  a26533a );
 a26538a <=( A269  and  A266 );
 a26539a <=( (not A265)  and  a26538a );
 a26540a <=( a26539a  and  a26534a );
 a26543a <=( (not A167)  and  (not A169) );
 a26547a <=( A200  and  (not A199) );
 a26548a <=( (not A166)  and  a26547a );
 a26549a <=( a26548a  and  a26543a );
 a26553a <=( A234  and  A233 );
 a26554a <=( A203  and  a26553a );
 a26558a <=( A269  and  (not A266) );
 a26559a <=( A265  and  a26558a );
 a26560a <=( a26559a  and  a26554a );
 a26563a <=( (not A167)  and  (not A169) );
 a26567a <=( A200  and  (not A199) );
 a26568a <=( (not A166)  and  a26567a );
 a26569a <=( a26568a  and  a26563a );
 a26573a <=( A233  and  (not A232) );
 a26574a <=( A203  and  a26573a );
 a26578a <=( A300  and  A299 );
 a26579a <=( A236  and  a26578a );
 a26580a <=( a26579a  and  a26574a );
 a26583a <=( (not A167)  and  (not A169) );
 a26587a <=( A200  and  (not A199) );
 a26588a <=( (not A166)  and  a26587a );
 a26589a <=( a26588a  and  a26583a );
 a26593a <=( A233  and  (not A232) );
 a26594a <=( A203  and  a26593a );
 a26598a <=( A300  and  A298 );
 a26599a <=( A236  and  a26598a );
 a26600a <=( a26599a  and  a26594a );
 a26603a <=( (not A167)  and  (not A169) );
 a26607a <=( A200  and  (not A199) );
 a26608a <=( (not A166)  and  a26607a );
 a26609a <=( a26608a  and  a26603a );
 a26613a <=( A233  and  (not A232) );
 a26614a <=( A203  and  a26613a );
 a26618a <=( A267  and  A265 );
 a26619a <=( A236  and  a26618a );
 a26620a <=( a26619a  and  a26614a );
 a26623a <=( (not A167)  and  (not A169) );
 a26627a <=( A200  and  (not A199) );
 a26628a <=( (not A166)  and  a26627a );
 a26629a <=( a26628a  and  a26623a );
 a26633a <=( A233  and  (not A232) );
 a26634a <=( A203  and  a26633a );
 a26638a <=( A267  and  A266 );
 a26639a <=( A236  and  a26638a );
 a26640a <=( a26639a  and  a26634a );
 a26643a <=( (not A167)  and  (not A169) );
 a26647a <=( A200  and  (not A199) );
 a26648a <=( (not A166)  and  a26647a );
 a26649a <=( a26648a  and  a26643a );
 a26653a <=( (not A233)  and  A232 );
 a26654a <=( A203  and  a26653a );
 a26658a <=( A300  and  A299 );
 a26659a <=( A236  and  a26658a );
 a26660a <=( a26659a  and  a26654a );
 a26663a <=( (not A167)  and  (not A169) );
 a26667a <=( A200  and  (not A199) );
 a26668a <=( (not A166)  and  a26667a );
 a26669a <=( a26668a  and  a26663a );
 a26673a <=( (not A233)  and  A232 );
 a26674a <=( A203  and  a26673a );
 a26678a <=( A300  and  A298 );
 a26679a <=( A236  and  a26678a );
 a26680a <=( a26679a  and  a26674a );
 a26683a <=( (not A167)  and  (not A169) );
 a26687a <=( A200  and  (not A199) );
 a26688a <=( (not A166)  and  a26687a );
 a26689a <=( a26688a  and  a26683a );
 a26693a <=( (not A233)  and  A232 );
 a26694a <=( A203  and  a26693a );
 a26698a <=( A267  and  A265 );
 a26699a <=( A236  and  a26698a );
 a26700a <=( a26699a  and  a26694a );
 a26703a <=( (not A167)  and  (not A169) );
 a26707a <=( A200  and  (not A199) );
 a26708a <=( (not A166)  and  a26707a );
 a26709a <=( a26708a  and  a26703a );
 a26713a <=( (not A233)  and  A232 );
 a26714a <=( A203  and  a26713a );
 a26718a <=( A267  and  A266 );
 a26719a <=( A236  and  a26718a );
 a26720a <=( a26719a  and  a26714a );
 a26723a <=( (not A167)  and  (not A169) );
 a26727a <=( (not A200)  and  A199 );
 a26728a <=( (not A166)  and  a26727a );
 a26729a <=( a26728a  and  a26723a );
 a26733a <=( A234  and  A232 );
 a26734a <=( A203  and  a26733a );
 a26738a <=( A302  and  (not A299) );
 a26739a <=( A298  and  a26738a );
 a26740a <=( a26739a  and  a26734a );
 a26743a <=( (not A167)  and  (not A169) );
 a26747a <=( (not A200)  and  A199 );
 a26748a <=( (not A166)  and  a26747a );
 a26749a <=( a26748a  and  a26743a );
 a26753a <=( A234  and  A232 );
 a26754a <=( A203  and  a26753a );
 a26758a <=( A302  and  A299 );
 a26759a <=( (not A298)  and  a26758a );
 a26760a <=( a26759a  and  a26754a );
 a26763a <=( (not A167)  and  (not A169) );
 a26767a <=( (not A200)  and  A199 );
 a26768a <=( (not A166)  and  a26767a );
 a26769a <=( a26768a  and  a26763a );
 a26773a <=( A234  and  A232 );
 a26774a <=( A203  and  a26773a );
 a26778a <=( A269  and  A266 );
 a26779a <=( (not A265)  and  a26778a );
 a26780a <=( a26779a  and  a26774a );
 a26783a <=( (not A167)  and  (not A169) );
 a26787a <=( (not A200)  and  A199 );
 a26788a <=( (not A166)  and  a26787a );
 a26789a <=( a26788a  and  a26783a );
 a26793a <=( A234  and  A232 );
 a26794a <=( A203  and  a26793a );
 a26798a <=( A269  and  (not A266) );
 a26799a <=( A265  and  a26798a );
 a26800a <=( a26799a  and  a26794a );
 a26803a <=( (not A167)  and  (not A169) );
 a26807a <=( (not A200)  and  A199 );
 a26808a <=( (not A166)  and  a26807a );
 a26809a <=( a26808a  and  a26803a );
 a26813a <=( A234  and  A233 );
 a26814a <=( A203  and  a26813a );
 a26818a <=( A302  and  (not A299) );
 a26819a <=( A298  and  a26818a );
 a26820a <=( a26819a  and  a26814a );
 a26823a <=( (not A167)  and  (not A169) );
 a26827a <=( (not A200)  and  A199 );
 a26828a <=( (not A166)  and  a26827a );
 a26829a <=( a26828a  and  a26823a );
 a26833a <=( A234  and  A233 );
 a26834a <=( A203  and  a26833a );
 a26838a <=( A302  and  A299 );
 a26839a <=( (not A298)  and  a26838a );
 a26840a <=( a26839a  and  a26834a );
 a26843a <=( (not A167)  and  (not A169) );
 a26847a <=( (not A200)  and  A199 );
 a26848a <=( (not A166)  and  a26847a );
 a26849a <=( a26848a  and  a26843a );
 a26853a <=( A234  and  A233 );
 a26854a <=( A203  and  a26853a );
 a26858a <=( A269  and  A266 );
 a26859a <=( (not A265)  and  a26858a );
 a26860a <=( a26859a  and  a26854a );
 a26863a <=( (not A167)  and  (not A169) );
 a26867a <=( (not A200)  and  A199 );
 a26868a <=( (not A166)  and  a26867a );
 a26869a <=( a26868a  and  a26863a );
 a26873a <=( A234  and  A233 );
 a26874a <=( A203  and  a26873a );
 a26878a <=( A269  and  (not A266) );
 a26879a <=( A265  and  a26878a );
 a26880a <=( a26879a  and  a26874a );
 a26883a <=( (not A167)  and  (not A169) );
 a26887a <=( (not A200)  and  A199 );
 a26888a <=( (not A166)  and  a26887a );
 a26889a <=( a26888a  and  a26883a );
 a26893a <=( A233  and  (not A232) );
 a26894a <=( A203  and  a26893a );
 a26898a <=( A300  and  A299 );
 a26899a <=( A236  and  a26898a );
 a26900a <=( a26899a  and  a26894a );
 a26903a <=( (not A167)  and  (not A169) );
 a26907a <=( (not A200)  and  A199 );
 a26908a <=( (not A166)  and  a26907a );
 a26909a <=( a26908a  and  a26903a );
 a26913a <=( A233  and  (not A232) );
 a26914a <=( A203  and  a26913a );
 a26918a <=( A300  and  A298 );
 a26919a <=( A236  and  a26918a );
 a26920a <=( a26919a  and  a26914a );
 a26923a <=( (not A167)  and  (not A169) );
 a26927a <=( (not A200)  and  A199 );
 a26928a <=( (not A166)  and  a26927a );
 a26929a <=( a26928a  and  a26923a );
 a26933a <=( A233  and  (not A232) );
 a26934a <=( A203  and  a26933a );
 a26938a <=( A267  and  A265 );
 a26939a <=( A236  and  a26938a );
 a26940a <=( a26939a  and  a26934a );
 a26943a <=( (not A167)  and  (not A169) );
 a26947a <=( (not A200)  and  A199 );
 a26948a <=( (not A166)  and  a26947a );
 a26949a <=( a26948a  and  a26943a );
 a26953a <=( A233  and  (not A232) );
 a26954a <=( A203  and  a26953a );
 a26958a <=( A267  and  A266 );
 a26959a <=( A236  and  a26958a );
 a26960a <=( a26959a  and  a26954a );
 a26963a <=( (not A167)  and  (not A169) );
 a26967a <=( (not A200)  and  A199 );
 a26968a <=( (not A166)  and  a26967a );
 a26969a <=( a26968a  and  a26963a );
 a26973a <=( (not A233)  and  A232 );
 a26974a <=( A203  and  a26973a );
 a26978a <=( A300  and  A299 );
 a26979a <=( A236  and  a26978a );
 a26980a <=( a26979a  and  a26974a );
 a26983a <=( (not A167)  and  (not A169) );
 a26987a <=( (not A200)  and  A199 );
 a26988a <=( (not A166)  and  a26987a );
 a26989a <=( a26988a  and  a26983a );
 a26993a <=( (not A233)  and  A232 );
 a26994a <=( A203  and  a26993a );
 a26998a <=( A300  and  A298 );
 a26999a <=( A236  and  a26998a );
 a27000a <=( a26999a  and  a26994a );
 a27003a <=( (not A167)  and  (not A169) );
 a27007a <=( (not A200)  and  A199 );
 a27008a <=( (not A166)  and  a27007a );
 a27009a <=( a27008a  and  a27003a );
 a27013a <=( (not A233)  and  A232 );
 a27014a <=( A203  and  a27013a );
 a27018a <=( A267  and  A265 );
 a27019a <=( A236  and  a27018a );
 a27020a <=( a27019a  and  a27014a );
 a27023a <=( (not A167)  and  (not A169) );
 a27027a <=( (not A200)  and  A199 );
 a27028a <=( (not A166)  and  a27027a );
 a27029a <=( a27028a  and  a27023a );
 a27033a <=( (not A233)  and  A232 );
 a27034a <=( A203  and  a27033a );
 a27038a <=( A267  and  A266 );
 a27039a <=( A236  and  a27038a );
 a27040a <=( a27039a  and  a27034a );
 a27043a <=( (not A168)  and  (not A169) );
 a27047a <=( A202  and  A166 );
 a27048a <=( A167  and  a27047a );
 a27049a <=( a27048a  and  a27043a );
 a27053a <=( A236  and  A233 );
 a27054a <=( (not A232)  and  a27053a );
 a27058a <=( A302  and  (not A299) );
 a27059a <=( A298  and  a27058a );
 a27060a <=( a27059a  and  a27054a );
 a27063a <=( (not A168)  and  (not A169) );
 a27067a <=( A202  and  A166 );
 a27068a <=( A167  and  a27067a );
 a27069a <=( a27068a  and  a27063a );
 a27073a <=( A236  and  A233 );
 a27074a <=( (not A232)  and  a27073a );
 a27078a <=( A302  and  A299 );
 a27079a <=( (not A298)  and  a27078a );
 a27080a <=( a27079a  and  a27074a );
 a27083a <=( (not A168)  and  (not A169) );
 a27087a <=( A202  and  A166 );
 a27088a <=( A167  and  a27087a );
 a27089a <=( a27088a  and  a27083a );
 a27093a <=( A236  and  A233 );
 a27094a <=( (not A232)  and  a27093a );
 a27098a <=( A269  and  A266 );
 a27099a <=( (not A265)  and  a27098a );
 a27100a <=( a27099a  and  a27094a );
 a27103a <=( (not A168)  and  (not A169) );
 a27107a <=( A202  and  A166 );
 a27108a <=( A167  and  a27107a );
 a27109a <=( a27108a  and  a27103a );
 a27113a <=( A236  and  A233 );
 a27114a <=( (not A232)  and  a27113a );
 a27118a <=( A269  and  (not A266) );
 a27119a <=( A265  and  a27118a );
 a27120a <=( a27119a  and  a27114a );
 a27123a <=( (not A168)  and  (not A169) );
 a27127a <=( A202  and  A166 );
 a27128a <=( A167  and  a27127a );
 a27129a <=( a27128a  and  a27123a );
 a27133a <=( A236  and  (not A233) );
 a27134a <=( A232  and  a27133a );
 a27138a <=( A302  and  (not A299) );
 a27139a <=( A298  and  a27138a );
 a27140a <=( a27139a  and  a27134a );
 a27143a <=( (not A168)  and  (not A169) );
 a27147a <=( A202  and  A166 );
 a27148a <=( A167  and  a27147a );
 a27149a <=( a27148a  and  a27143a );
 a27153a <=( A236  and  (not A233) );
 a27154a <=( A232  and  a27153a );
 a27158a <=( A302  and  A299 );
 a27159a <=( (not A298)  and  a27158a );
 a27160a <=( a27159a  and  a27154a );
 a27163a <=( (not A168)  and  (not A169) );
 a27167a <=( A202  and  A166 );
 a27168a <=( A167  and  a27167a );
 a27169a <=( a27168a  and  a27163a );
 a27173a <=( A236  and  (not A233) );
 a27174a <=( A232  and  a27173a );
 a27178a <=( A269  and  A266 );
 a27179a <=( (not A265)  and  a27178a );
 a27180a <=( a27179a  and  a27174a );
 a27183a <=( (not A168)  and  (not A169) );
 a27187a <=( A202  and  A166 );
 a27188a <=( A167  and  a27187a );
 a27189a <=( a27188a  and  a27183a );
 a27193a <=( A236  and  (not A233) );
 a27194a <=( A232  and  a27193a );
 a27198a <=( A269  and  (not A266) );
 a27199a <=( A265  and  a27198a );
 a27200a <=( a27199a  and  a27194a );
 a27203a <=( (not A168)  and  (not A169) );
 a27207a <=( A199  and  A166 );
 a27208a <=( A167  and  a27207a );
 a27209a <=( a27208a  and  a27203a );
 a27213a <=( A234  and  A232 );
 a27214a <=( A201  and  a27213a );
 a27218a <=( A302  and  (not A299) );
 a27219a <=( A298  and  a27218a );
 a27220a <=( a27219a  and  a27214a );
 a27223a <=( (not A168)  and  (not A169) );
 a27227a <=( A199  and  A166 );
 a27228a <=( A167  and  a27227a );
 a27229a <=( a27228a  and  a27223a );
 a27233a <=( A234  and  A232 );
 a27234a <=( A201  and  a27233a );
 a27238a <=( A302  and  A299 );
 a27239a <=( (not A298)  and  a27238a );
 a27240a <=( a27239a  and  a27234a );
 a27243a <=( (not A168)  and  (not A169) );
 a27247a <=( A199  and  A166 );
 a27248a <=( A167  and  a27247a );
 a27249a <=( a27248a  and  a27243a );
 a27253a <=( A234  and  A232 );
 a27254a <=( A201  and  a27253a );
 a27258a <=( A269  and  A266 );
 a27259a <=( (not A265)  and  a27258a );
 a27260a <=( a27259a  and  a27254a );
 a27263a <=( (not A168)  and  (not A169) );
 a27267a <=( A199  and  A166 );
 a27268a <=( A167  and  a27267a );
 a27269a <=( a27268a  and  a27263a );
 a27273a <=( A234  and  A232 );
 a27274a <=( A201  and  a27273a );
 a27278a <=( A269  and  (not A266) );
 a27279a <=( A265  and  a27278a );
 a27280a <=( a27279a  and  a27274a );
 a27283a <=( (not A168)  and  (not A169) );
 a27287a <=( A199  and  A166 );
 a27288a <=( A167  and  a27287a );
 a27289a <=( a27288a  and  a27283a );
 a27293a <=( A234  and  A233 );
 a27294a <=( A201  and  a27293a );
 a27298a <=( A302  and  (not A299) );
 a27299a <=( A298  and  a27298a );
 a27300a <=( a27299a  and  a27294a );
 a27303a <=( (not A168)  and  (not A169) );
 a27307a <=( A199  and  A166 );
 a27308a <=( A167  and  a27307a );
 a27309a <=( a27308a  and  a27303a );
 a27313a <=( A234  and  A233 );
 a27314a <=( A201  and  a27313a );
 a27318a <=( A302  and  A299 );
 a27319a <=( (not A298)  and  a27318a );
 a27320a <=( a27319a  and  a27314a );
 a27323a <=( (not A168)  and  (not A169) );
 a27327a <=( A199  and  A166 );
 a27328a <=( A167  and  a27327a );
 a27329a <=( a27328a  and  a27323a );
 a27333a <=( A234  and  A233 );
 a27334a <=( A201  and  a27333a );
 a27338a <=( A269  and  A266 );
 a27339a <=( (not A265)  and  a27338a );
 a27340a <=( a27339a  and  a27334a );
 a27343a <=( (not A168)  and  (not A169) );
 a27347a <=( A199  and  A166 );
 a27348a <=( A167  and  a27347a );
 a27349a <=( a27348a  and  a27343a );
 a27353a <=( A234  and  A233 );
 a27354a <=( A201  and  a27353a );
 a27358a <=( A269  and  (not A266) );
 a27359a <=( A265  and  a27358a );
 a27360a <=( a27359a  and  a27354a );
 a27363a <=( (not A168)  and  (not A169) );
 a27367a <=( A199  and  A166 );
 a27368a <=( A167  and  a27367a );
 a27369a <=( a27368a  and  a27363a );
 a27373a <=( A233  and  (not A232) );
 a27374a <=( A201  and  a27373a );
 a27378a <=( A300  and  A299 );
 a27379a <=( A236  and  a27378a );
 a27380a <=( a27379a  and  a27374a );
 a27383a <=( (not A168)  and  (not A169) );
 a27387a <=( A199  and  A166 );
 a27388a <=( A167  and  a27387a );
 a27389a <=( a27388a  and  a27383a );
 a27393a <=( A233  and  (not A232) );
 a27394a <=( A201  and  a27393a );
 a27398a <=( A300  and  A298 );
 a27399a <=( A236  and  a27398a );
 a27400a <=( a27399a  and  a27394a );
 a27403a <=( (not A168)  and  (not A169) );
 a27407a <=( A199  and  A166 );
 a27408a <=( A167  and  a27407a );
 a27409a <=( a27408a  and  a27403a );
 a27413a <=( A233  and  (not A232) );
 a27414a <=( A201  and  a27413a );
 a27418a <=( A267  and  A265 );
 a27419a <=( A236  and  a27418a );
 a27420a <=( a27419a  and  a27414a );
 a27423a <=( (not A168)  and  (not A169) );
 a27427a <=( A199  and  A166 );
 a27428a <=( A167  and  a27427a );
 a27429a <=( a27428a  and  a27423a );
 a27433a <=( A233  and  (not A232) );
 a27434a <=( A201  and  a27433a );
 a27438a <=( A267  and  A266 );
 a27439a <=( A236  and  a27438a );
 a27440a <=( a27439a  and  a27434a );
 a27443a <=( (not A168)  and  (not A169) );
 a27447a <=( A199  and  A166 );
 a27448a <=( A167  and  a27447a );
 a27449a <=( a27448a  and  a27443a );
 a27453a <=( (not A233)  and  A232 );
 a27454a <=( A201  and  a27453a );
 a27458a <=( A300  and  A299 );
 a27459a <=( A236  and  a27458a );
 a27460a <=( a27459a  and  a27454a );
 a27463a <=( (not A168)  and  (not A169) );
 a27467a <=( A199  and  A166 );
 a27468a <=( A167  and  a27467a );
 a27469a <=( a27468a  and  a27463a );
 a27473a <=( (not A233)  and  A232 );
 a27474a <=( A201  and  a27473a );
 a27478a <=( A300  and  A298 );
 a27479a <=( A236  and  a27478a );
 a27480a <=( a27479a  and  a27474a );
 a27483a <=( (not A168)  and  (not A169) );
 a27487a <=( A199  and  A166 );
 a27488a <=( A167  and  a27487a );
 a27489a <=( a27488a  and  a27483a );
 a27493a <=( (not A233)  and  A232 );
 a27494a <=( A201  and  a27493a );
 a27498a <=( A267  and  A265 );
 a27499a <=( A236  and  a27498a );
 a27500a <=( a27499a  and  a27494a );
 a27503a <=( (not A168)  and  (not A169) );
 a27507a <=( A199  and  A166 );
 a27508a <=( A167  and  a27507a );
 a27509a <=( a27508a  and  a27503a );
 a27513a <=( (not A233)  and  A232 );
 a27514a <=( A201  and  a27513a );
 a27518a <=( A267  and  A266 );
 a27519a <=( A236  and  a27518a );
 a27520a <=( a27519a  and  a27514a );
 a27523a <=( (not A168)  and  (not A169) );
 a27527a <=( A200  and  A166 );
 a27528a <=( A167  and  a27527a );
 a27529a <=( a27528a  and  a27523a );
 a27533a <=( A234  and  A232 );
 a27534a <=( A201  and  a27533a );
 a27538a <=( A302  and  (not A299) );
 a27539a <=( A298  and  a27538a );
 a27540a <=( a27539a  and  a27534a );
 a27543a <=( (not A168)  and  (not A169) );
 a27547a <=( A200  and  A166 );
 a27548a <=( A167  and  a27547a );
 a27549a <=( a27548a  and  a27543a );
 a27553a <=( A234  and  A232 );
 a27554a <=( A201  and  a27553a );
 a27558a <=( A302  and  A299 );
 a27559a <=( (not A298)  and  a27558a );
 a27560a <=( a27559a  and  a27554a );
 a27563a <=( (not A168)  and  (not A169) );
 a27567a <=( A200  and  A166 );
 a27568a <=( A167  and  a27567a );
 a27569a <=( a27568a  and  a27563a );
 a27573a <=( A234  and  A232 );
 a27574a <=( A201  and  a27573a );
 a27578a <=( A269  and  A266 );
 a27579a <=( (not A265)  and  a27578a );
 a27580a <=( a27579a  and  a27574a );
 a27583a <=( (not A168)  and  (not A169) );
 a27587a <=( A200  and  A166 );
 a27588a <=( A167  and  a27587a );
 a27589a <=( a27588a  and  a27583a );
 a27593a <=( A234  and  A232 );
 a27594a <=( A201  and  a27593a );
 a27598a <=( A269  and  (not A266) );
 a27599a <=( A265  and  a27598a );
 a27600a <=( a27599a  and  a27594a );
 a27603a <=( (not A168)  and  (not A169) );
 a27607a <=( A200  and  A166 );
 a27608a <=( A167  and  a27607a );
 a27609a <=( a27608a  and  a27603a );
 a27613a <=( A234  and  A233 );
 a27614a <=( A201  and  a27613a );
 a27618a <=( A302  and  (not A299) );
 a27619a <=( A298  and  a27618a );
 a27620a <=( a27619a  and  a27614a );
 a27623a <=( (not A168)  and  (not A169) );
 a27627a <=( A200  and  A166 );
 a27628a <=( A167  and  a27627a );
 a27629a <=( a27628a  and  a27623a );
 a27633a <=( A234  and  A233 );
 a27634a <=( A201  and  a27633a );
 a27638a <=( A302  and  A299 );
 a27639a <=( (not A298)  and  a27638a );
 a27640a <=( a27639a  and  a27634a );
 a27643a <=( (not A168)  and  (not A169) );
 a27647a <=( A200  and  A166 );
 a27648a <=( A167  and  a27647a );
 a27649a <=( a27648a  and  a27643a );
 a27653a <=( A234  and  A233 );
 a27654a <=( A201  and  a27653a );
 a27658a <=( A269  and  A266 );
 a27659a <=( (not A265)  and  a27658a );
 a27660a <=( a27659a  and  a27654a );
 a27663a <=( (not A168)  and  (not A169) );
 a27667a <=( A200  and  A166 );
 a27668a <=( A167  and  a27667a );
 a27669a <=( a27668a  and  a27663a );
 a27673a <=( A234  and  A233 );
 a27674a <=( A201  and  a27673a );
 a27678a <=( A269  and  (not A266) );
 a27679a <=( A265  and  a27678a );
 a27680a <=( a27679a  and  a27674a );
 a27683a <=( (not A168)  and  (not A169) );
 a27687a <=( A200  and  A166 );
 a27688a <=( A167  and  a27687a );
 a27689a <=( a27688a  and  a27683a );
 a27693a <=( A233  and  (not A232) );
 a27694a <=( A201  and  a27693a );
 a27698a <=( A300  and  A299 );
 a27699a <=( A236  and  a27698a );
 a27700a <=( a27699a  and  a27694a );
 a27703a <=( (not A168)  and  (not A169) );
 a27707a <=( A200  and  A166 );
 a27708a <=( A167  and  a27707a );
 a27709a <=( a27708a  and  a27703a );
 a27713a <=( A233  and  (not A232) );
 a27714a <=( A201  and  a27713a );
 a27718a <=( A300  and  A298 );
 a27719a <=( A236  and  a27718a );
 a27720a <=( a27719a  and  a27714a );
 a27723a <=( (not A168)  and  (not A169) );
 a27727a <=( A200  and  A166 );
 a27728a <=( A167  and  a27727a );
 a27729a <=( a27728a  and  a27723a );
 a27733a <=( A233  and  (not A232) );
 a27734a <=( A201  and  a27733a );
 a27738a <=( A267  and  A265 );
 a27739a <=( A236  and  a27738a );
 a27740a <=( a27739a  and  a27734a );
 a27743a <=( (not A168)  and  (not A169) );
 a27747a <=( A200  and  A166 );
 a27748a <=( A167  and  a27747a );
 a27749a <=( a27748a  and  a27743a );
 a27753a <=( A233  and  (not A232) );
 a27754a <=( A201  and  a27753a );
 a27758a <=( A267  and  A266 );
 a27759a <=( A236  and  a27758a );
 a27760a <=( a27759a  and  a27754a );
 a27763a <=( (not A168)  and  (not A169) );
 a27767a <=( A200  and  A166 );
 a27768a <=( A167  and  a27767a );
 a27769a <=( a27768a  and  a27763a );
 a27773a <=( (not A233)  and  A232 );
 a27774a <=( A201  and  a27773a );
 a27778a <=( A300  and  A299 );
 a27779a <=( A236  and  a27778a );
 a27780a <=( a27779a  and  a27774a );
 a27783a <=( (not A168)  and  (not A169) );
 a27787a <=( A200  and  A166 );
 a27788a <=( A167  and  a27787a );
 a27789a <=( a27788a  and  a27783a );
 a27793a <=( (not A233)  and  A232 );
 a27794a <=( A201  and  a27793a );
 a27798a <=( A300  and  A298 );
 a27799a <=( A236  and  a27798a );
 a27800a <=( a27799a  and  a27794a );
 a27803a <=( (not A168)  and  (not A169) );
 a27807a <=( A200  and  A166 );
 a27808a <=( A167  and  a27807a );
 a27809a <=( a27808a  and  a27803a );
 a27813a <=( (not A233)  and  A232 );
 a27814a <=( A201  and  a27813a );
 a27818a <=( A267  and  A265 );
 a27819a <=( A236  and  a27818a );
 a27820a <=( a27819a  and  a27814a );
 a27823a <=( (not A168)  and  (not A169) );
 a27827a <=( A200  and  A166 );
 a27828a <=( A167  and  a27827a );
 a27829a <=( a27828a  and  a27823a );
 a27833a <=( (not A233)  and  A232 );
 a27834a <=( A201  and  a27833a );
 a27838a <=( A267  and  A266 );
 a27839a <=( A236  and  a27838a );
 a27840a <=( a27839a  and  a27834a );
 a27843a <=( (not A168)  and  (not A169) );
 a27847a <=( (not A199)  and  A166 );
 a27848a <=( A167  and  a27847a );
 a27849a <=( a27848a  and  a27843a );
 a27853a <=( A235  and  A203 );
 a27854a <=( A200  and  a27853a );
 a27858a <=( A302  and  (not A299) );
 a27859a <=( A298  and  a27858a );
 a27860a <=( a27859a  and  a27854a );
 a27863a <=( (not A168)  and  (not A169) );
 a27867a <=( (not A199)  and  A166 );
 a27868a <=( A167  and  a27867a );
 a27869a <=( a27868a  and  a27863a );
 a27873a <=( A235  and  A203 );
 a27874a <=( A200  and  a27873a );
 a27878a <=( A302  and  A299 );
 a27879a <=( (not A298)  and  a27878a );
 a27880a <=( a27879a  and  a27874a );
 a27883a <=( (not A168)  and  (not A169) );
 a27887a <=( (not A199)  and  A166 );
 a27888a <=( A167  and  a27887a );
 a27889a <=( a27888a  and  a27883a );
 a27893a <=( A235  and  A203 );
 a27894a <=( A200  and  a27893a );
 a27898a <=( A269  and  A266 );
 a27899a <=( (not A265)  and  a27898a );
 a27900a <=( a27899a  and  a27894a );
 a27903a <=( (not A168)  and  (not A169) );
 a27907a <=( (not A199)  and  A166 );
 a27908a <=( A167  and  a27907a );
 a27909a <=( a27908a  and  a27903a );
 a27913a <=( A235  and  A203 );
 a27914a <=( A200  and  a27913a );
 a27918a <=( A269  and  (not A266) );
 a27919a <=( A265  and  a27918a );
 a27920a <=( a27919a  and  a27914a );
 a27923a <=( (not A168)  and  (not A169) );
 a27927a <=( (not A199)  and  A166 );
 a27928a <=( A167  and  a27927a );
 a27929a <=( a27928a  and  a27923a );
 a27933a <=( A232  and  A203 );
 a27934a <=( A200  and  a27933a );
 a27938a <=( A300  and  A299 );
 a27939a <=( A234  and  a27938a );
 a27940a <=( a27939a  and  a27934a );
 a27943a <=( (not A168)  and  (not A169) );
 a27947a <=( (not A199)  and  A166 );
 a27948a <=( A167  and  a27947a );
 a27949a <=( a27948a  and  a27943a );
 a27953a <=( A232  and  A203 );
 a27954a <=( A200  and  a27953a );
 a27958a <=( A300  and  A298 );
 a27959a <=( A234  and  a27958a );
 a27960a <=( a27959a  and  a27954a );
 a27963a <=( (not A168)  and  (not A169) );
 a27967a <=( (not A199)  and  A166 );
 a27968a <=( A167  and  a27967a );
 a27969a <=( a27968a  and  a27963a );
 a27973a <=( A232  and  A203 );
 a27974a <=( A200  and  a27973a );
 a27978a <=( A267  and  A265 );
 a27979a <=( A234  and  a27978a );
 a27980a <=( a27979a  and  a27974a );
 a27983a <=( (not A168)  and  (not A169) );
 a27987a <=( (not A199)  and  A166 );
 a27988a <=( A167  and  a27987a );
 a27989a <=( a27988a  and  a27983a );
 a27993a <=( A232  and  A203 );
 a27994a <=( A200  and  a27993a );
 a27998a <=( A267  and  A266 );
 a27999a <=( A234  and  a27998a );
 a28000a <=( a27999a  and  a27994a );
 a28003a <=( (not A168)  and  (not A169) );
 a28007a <=( (not A199)  and  A166 );
 a28008a <=( A167  and  a28007a );
 a28009a <=( a28008a  and  a28003a );
 a28013a <=( A233  and  A203 );
 a28014a <=( A200  and  a28013a );
 a28018a <=( A300  and  A299 );
 a28019a <=( A234  and  a28018a );
 a28020a <=( a28019a  and  a28014a );
 a28023a <=( (not A168)  and  (not A169) );
 a28027a <=( (not A199)  and  A166 );
 a28028a <=( A167  and  a28027a );
 a28029a <=( a28028a  and  a28023a );
 a28033a <=( A233  and  A203 );
 a28034a <=( A200  and  a28033a );
 a28038a <=( A300  and  A298 );
 a28039a <=( A234  and  a28038a );
 a28040a <=( a28039a  and  a28034a );
 a28043a <=( (not A168)  and  (not A169) );
 a28047a <=( (not A199)  and  A166 );
 a28048a <=( A167  and  a28047a );
 a28049a <=( a28048a  and  a28043a );
 a28053a <=( A233  and  A203 );
 a28054a <=( A200  and  a28053a );
 a28058a <=( A267  and  A265 );
 a28059a <=( A234  and  a28058a );
 a28060a <=( a28059a  and  a28054a );
 a28063a <=( (not A168)  and  (not A169) );
 a28067a <=( (not A199)  and  A166 );
 a28068a <=( A167  and  a28067a );
 a28069a <=( a28068a  and  a28063a );
 a28073a <=( A233  and  A203 );
 a28074a <=( A200  and  a28073a );
 a28078a <=( A267  and  A266 );
 a28079a <=( A234  and  a28078a );
 a28080a <=( a28079a  and  a28074a );
 a28083a <=( (not A168)  and  (not A169) );
 a28087a <=( (not A199)  and  A166 );
 a28088a <=( A167  and  a28087a );
 a28089a <=( a28088a  and  a28083a );
 a28093a <=( (not A232)  and  A203 );
 a28094a <=( A200  and  a28093a );
 a28098a <=( A301  and  A236 );
 a28099a <=( A233  and  a28098a );
 a28100a <=( a28099a  and  a28094a );
 a28103a <=( (not A168)  and  (not A169) );
 a28107a <=( (not A199)  and  A166 );
 a28108a <=( A167  and  a28107a );
 a28109a <=( a28108a  and  a28103a );
 a28113a <=( (not A232)  and  A203 );
 a28114a <=( A200  and  a28113a );
 a28118a <=( A268  and  A236 );
 a28119a <=( A233  and  a28118a );
 a28120a <=( a28119a  and  a28114a );
 a28123a <=( (not A168)  and  (not A169) );
 a28127a <=( (not A199)  and  A166 );
 a28128a <=( A167  and  a28127a );
 a28129a <=( a28128a  and  a28123a );
 a28133a <=( A232  and  A203 );
 a28134a <=( A200  and  a28133a );
 a28138a <=( A301  and  A236 );
 a28139a <=( (not A233)  and  a28138a );
 a28140a <=( a28139a  and  a28134a );
 a28143a <=( (not A168)  and  (not A169) );
 a28147a <=( (not A199)  and  A166 );
 a28148a <=( A167  and  a28147a );
 a28149a <=( a28148a  and  a28143a );
 a28153a <=( A232  and  A203 );
 a28154a <=( A200  and  a28153a );
 a28158a <=( A268  and  A236 );
 a28159a <=( (not A233)  and  a28158a );
 a28160a <=( a28159a  and  a28154a );
 a28163a <=( (not A168)  and  (not A169) );
 a28167a <=( A199  and  A166 );
 a28168a <=( A167  and  a28167a );
 a28169a <=( a28168a  and  a28163a );
 a28173a <=( A235  and  A203 );
 a28174a <=( (not A200)  and  a28173a );
 a28178a <=( A302  and  (not A299) );
 a28179a <=( A298  and  a28178a );
 a28180a <=( a28179a  and  a28174a );
 a28183a <=( (not A168)  and  (not A169) );
 a28187a <=( A199  and  A166 );
 a28188a <=( A167  and  a28187a );
 a28189a <=( a28188a  and  a28183a );
 a28193a <=( A235  and  A203 );
 a28194a <=( (not A200)  and  a28193a );
 a28198a <=( A302  and  A299 );
 a28199a <=( (not A298)  and  a28198a );
 a28200a <=( a28199a  and  a28194a );
 a28203a <=( (not A168)  and  (not A169) );
 a28207a <=( A199  and  A166 );
 a28208a <=( A167  and  a28207a );
 a28209a <=( a28208a  and  a28203a );
 a28213a <=( A235  and  A203 );
 a28214a <=( (not A200)  and  a28213a );
 a28218a <=( A269  and  A266 );
 a28219a <=( (not A265)  and  a28218a );
 a28220a <=( a28219a  and  a28214a );
 a28223a <=( (not A168)  and  (not A169) );
 a28227a <=( A199  and  A166 );
 a28228a <=( A167  and  a28227a );
 a28229a <=( a28228a  and  a28223a );
 a28233a <=( A235  and  A203 );
 a28234a <=( (not A200)  and  a28233a );
 a28238a <=( A269  and  (not A266) );
 a28239a <=( A265  and  a28238a );
 a28240a <=( a28239a  and  a28234a );
 a28243a <=( (not A168)  and  (not A169) );
 a28247a <=( A199  and  A166 );
 a28248a <=( A167  and  a28247a );
 a28249a <=( a28248a  and  a28243a );
 a28253a <=( A232  and  A203 );
 a28254a <=( (not A200)  and  a28253a );
 a28258a <=( A300  and  A299 );
 a28259a <=( A234  and  a28258a );
 a28260a <=( a28259a  and  a28254a );
 a28263a <=( (not A168)  and  (not A169) );
 a28267a <=( A199  and  A166 );
 a28268a <=( A167  and  a28267a );
 a28269a <=( a28268a  and  a28263a );
 a28273a <=( A232  and  A203 );
 a28274a <=( (not A200)  and  a28273a );
 a28278a <=( A300  and  A298 );
 a28279a <=( A234  and  a28278a );
 a28280a <=( a28279a  and  a28274a );
 a28283a <=( (not A168)  and  (not A169) );
 a28287a <=( A199  and  A166 );
 a28288a <=( A167  and  a28287a );
 a28289a <=( a28288a  and  a28283a );
 a28293a <=( A232  and  A203 );
 a28294a <=( (not A200)  and  a28293a );
 a28298a <=( A267  and  A265 );
 a28299a <=( A234  and  a28298a );
 a28300a <=( a28299a  and  a28294a );
 a28303a <=( (not A168)  and  (not A169) );
 a28307a <=( A199  and  A166 );
 a28308a <=( A167  and  a28307a );
 a28309a <=( a28308a  and  a28303a );
 a28313a <=( A232  and  A203 );
 a28314a <=( (not A200)  and  a28313a );
 a28318a <=( A267  and  A266 );
 a28319a <=( A234  and  a28318a );
 a28320a <=( a28319a  and  a28314a );
 a28323a <=( (not A168)  and  (not A169) );
 a28327a <=( A199  and  A166 );
 a28328a <=( A167  and  a28327a );
 a28329a <=( a28328a  and  a28323a );
 a28333a <=( A233  and  A203 );
 a28334a <=( (not A200)  and  a28333a );
 a28338a <=( A300  and  A299 );
 a28339a <=( A234  and  a28338a );
 a28340a <=( a28339a  and  a28334a );
 a28343a <=( (not A168)  and  (not A169) );
 a28347a <=( A199  and  A166 );
 a28348a <=( A167  and  a28347a );
 a28349a <=( a28348a  and  a28343a );
 a28353a <=( A233  and  A203 );
 a28354a <=( (not A200)  and  a28353a );
 a28358a <=( A300  and  A298 );
 a28359a <=( A234  and  a28358a );
 a28360a <=( a28359a  and  a28354a );
 a28363a <=( (not A168)  and  (not A169) );
 a28367a <=( A199  and  A166 );
 a28368a <=( A167  and  a28367a );
 a28369a <=( a28368a  and  a28363a );
 a28373a <=( A233  and  A203 );
 a28374a <=( (not A200)  and  a28373a );
 a28378a <=( A267  and  A265 );
 a28379a <=( A234  and  a28378a );
 a28380a <=( a28379a  and  a28374a );
 a28383a <=( (not A168)  and  (not A169) );
 a28387a <=( A199  and  A166 );
 a28388a <=( A167  and  a28387a );
 a28389a <=( a28388a  and  a28383a );
 a28393a <=( A233  and  A203 );
 a28394a <=( (not A200)  and  a28393a );
 a28398a <=( A267  and  A266 );
 a28399a <=( A234  and  a28398a );
 a28400a <=( a28399a  and  a28394a );
 a28403a <=( (not A168)  and  (not A169) );
 a28407a <=( A199  and  A166 );
 a28408a <=( A167  and  a28407a );
 a28409a <=( a28408a  and  a28403a );
 a28413a <=( (not A232)  and  A203 );
 a28414a <=( (not A200)  and  a28413a );
 a28418a <=( A301  and  A236 );
 a28419a <=( A233  and  a28418a );
 a28420a <=( a28419a  and  a28414a );
 a28423a <=( (not A168)  and  (not A169) );
 a28427a <=( A199  and  A166 );
 a28428a <=( A167  and  a28427a );
 a28429a <=( a28428a  and  a28423a );
 a28433a <=( (not A232)  and  A203 );
 a28434a <=( (not A200)  and  a28433a );
 a28438a <=( A268  and  A236 );
 a28439a <=( A233  and  a28438a );
 a28440a <=( a28439a  and  a28434a );
 a28443a <=( (not A168)  and  (not A169) );
 a28447a <=( A199  and  A166 );
 a28448a <=( A167  and  a28447a );
 a28449a <=( a28448a  and  a28443a );
 a28453a <=( A232  and  A203 );
 a28454a <=( (not A200)  and  a28453a );
 a28458a <=( A301  and  A236 );
 a28459a <=( (not A233)  and  a28458a );
 a28460a <=( a28459a  and  a28454a );
 a28463a <=( (not A168)  and  (not A169) );
 a28467a <=( A199  and  A166 );
 a28468a <=( A167  and  a28467a );
 a28469a <=( a28468a  and  a28463a );
 a28473a <=( A232  and  A203 );
 a28474a <=( (not A200)  and  a28473a );
 a28478a <=( A268  and  A236 );
 a28479a <=( (not A233)  and  a28478a );
 a28480a <=( a28479a  and  a28474a );
 a28483a <=( (not A169)  and  (not A170) );
 a28487a <=( A201  and  A199 );
 a28488a <=( (not A168)  and  a28487a );
 a28489a <=( a28488a  and  a28483a );
 a28493a <=( A236  and  A233 );
 a28494a <=( (not A232)  and  a28493a );
 a28498a <=( A302  and  (not A299) );
 a28499a <=( A298  and  a28498a );
 a28500a <=( a28499a  and  a28494a );
 a28503a <=( (not A169)  and  (not A170) );
 a28507a <=( A201  and  A199 );
 a28508a <=( (not A168)  and  a28507a );
 a28509a <=( a28508a  and  a28503a );
 a28513a <=( A236  and  A233 );
 a28514a <=( (not A232)  and  a28513a );
 a28518a <=( A302  and  A299 );
 a28519a <=( (not A298)  and  a28518a );
 a28520a <=( a28519a  and  a28514a );
 a28523a <=( (not A169)  and  (not A170) );
 a28527a <=( A201  and  A199 );
 a28528a <=( (not A168)  and  a28527a );
 a28529a <=( a28528a  and  a28523a );
 a28533a <=( A236  and  A233 );
 a28534a <=( (not A232)  and  a28533a );
 a28538a <=( A269  and  A266 );
 a28539a <=( (not A265)  and  a28538a );
 a28540a <=( a28539a  and  a28534a );
 a28543a <=( (not A169)  and  (not A170) );
 a28547a <=( A201  and  A199 );
 a28548a <=( (not A168)  and  a28547a );
 a28549a <=( a28548a  and  a28543a );
 a28553a <=( A236  and  A233 );
 a28554a <=( (not A232)  and  a28553a );
 a28558a <=( A269  and  (not A266) );
 a28559a <=( A265  and  a28558a );
 a28560a <=( a28559a  and  a28554a );
 a28563a <=( (not A169)  and  (not A170) );
 a28567a <=( A201  and  A199 );
 a28568a <=( (not A168)  and  a28567a );
 a28569a <=( a28568a  and  a28563a );
 a28573a <=( A236  and  (not A233) );
 a28574a <=( A232  and  a28573a );
 a28578a <=( A302  and  (not A299) );
 a28579a <=( A298  and  a28578a );
 a28580a <=( a28579a  and  a28574a );
 a28583a <=( (not A169)  and  (not A170) );
 a28587a <=( A201  and  A199 );
 a28588a <=( (not A168)  and  a28587a );
 a28589a <=( a28588a  and  a28583a );
 a28593a <=( A236  and  (not A233) );
 a28594a <=( A232  and  a28593a );
 a28598a <=( A302  and  A299 );
 a28599a <=( (not A298)  and  a28598a );
 a28600a <=( a28599a  and  a28594a );
 a28603a <=( (not A169)  and  (not A170) );
 a28607a <=( A201  and  A199 );
 a28608a <=( (not A168)  and  a28607a );
 a28609a <=( a28608a  and  a28603a );
 a28613a <=( A236  and  (not A233) );
 a28614a <=( A232  and  a28613a );
 a28618a <=( A269  and  A266 );
 a28619a <=( (not A265)  and  a28618a );
 a28620a <=( a28619a  and  a28614a );
 a28623a <=( (not A169)  and  (not A170) );
 a28627a <=( A201  and  A199 );
 a28628a <=( (not A168)  and  a28627a );
 a28629a <=( a28628a  and  a28623a );
 a28633a <=( A236  and  (not A233) );
 a28634a <=( A232  and  a28633a );
 a28638a <=( A269  and  (not A266) );
 a28639a <=( A265  and  a28638a );
 a28640a <=( a28639a  and  a28634a );
 a28643a <=( (not A169)  and  (not A170) );
 a28647a <=( A201  and  A200 );
 a28648a <=( (not A168)  and  a28647a );
 a28649a <=( a28648a  and  a28643a );
 a28653a <=( A236  and  A233 );
 a28654a <=( (not A232)  and  a28653a );
 a28658a <=( A302  and  (not A299) );
 a28659a <=( A298  and  a28658a );
 a28660a <=( a28659a  and  a28654a );
 a28663a <=( (not A169)  and  (not A170) );
 a28667a <=( A201  and  A200 );
 a28668a <=( (not A168)  and  a28667a );
 a28669a <=( a28668a  and  a28663a );
 a28673a <=( A236  and  A233 );
 a28674a <=( (not A232)  and  a28673a );
 a28678a <=( A302  and  A299 );
 a28679a <=( (not A298)  and  a28678a );
 a28680a <=( a28679a  and  a28674a );
 a28683a <=( (not A169)  and  (not A170) );
 a28687a <=( A201  and  A200 );
 a28688a <=( (not A168)  and  a28687a );
 a28689a <=( a28688a  and  a28683a );
 a28693a <=( A236  and  A233 );
 a28694a <=( (not A232)  and  a28693a );
 a28698a <=( A269  and  A266 );
 a28699a <=( (not A265)  and  a28698a );
 a28700a <=( a28699a  and  a28694a );
 a28703a <=( (not A169)  and  (not A170) );
 a28707a <=( A201  and  A200 );
 a28708a <=( (not A168)  and  a28707a );
 a28709a <=( a28708a  and  a28703a );
 a28713a <=( A236  and  A233 );
 a28714a <=( (not A232)  and  a28713a );
 a28718a <=( A269  and  (not A266) );
 a28719a <=( A265  and  a28718a );
 a28720a <=( a28719a  and  a28714a );
 a28723a <=( (not A169)  and  (not A170) );
 a28727a <=( A201  and  A200 );
 a28728a <=( (not A168)  and  a28727a );
 a28729a <=( a28728a  and  a28723a );
 a28733a <=( A236  and  (not A233) );
 a28734a <=( A232  and  a28733a );
 a28738a <=( A302  and  (not A299) );
 a28739a <=( A298  and  a28738a );
 a28740a <=( a28739a  and  a28734a );
 a28743a <=( (not A169)  and  (not A170) );
 a28747a <=( A201  and  A200 );
 a28748a <=( (not A168)  and  a28747a );
 a28749a <=( a28748a  and  a28743a );
 a28753a <=( A236  and  (not A233) );
 a28754a <=( A232  and  a28753a );
 a28758a <=( A302  and  A299 );
 a28759a <=( (not A298)  and  a28758a );
 a28760a <=( a28759a  and  a28754a );
 a28763a <=( (not A169)  and  (not A170) );
 a28767a <=( A201  and  A200 );
 a28768a <=( (not A168)  and  a28767a );
 a28769a <=( a28768a  and  a28763a );
 a28773a <=( A236  and  (not A233) );
 a28774a <=( A232  and  a28773a );
 a28778a <=( A269  and  A266 );
 a28779a <=( (not A265)  and  a28778a );
 a28780a <=( a28779a  and  a28774a );
 a28783a <=( (not A169)  and  (not A170) );
 a28787a <=( A201  and  A200 );
 a28788a <=( (not A168)  and  a28787a );
 a28789a <=( a28788a  and  a28783a );
 a28793a <=( A236  and  (not A233) );
 a28794a <=( A232  and  a28793a );
 a28798a <=( A269  and  (not A266) );
 a28799a <=( A265  and  a28798a );
 a28800a <=( a28799a  and  a28794a );
 a28803a <=( (not A169)  and  (not A170) );
 a28807a <=( A200  and  (not A199) );
 a28808a <=( (not A168)  and  a28807a );
 a28809a <=( a28808a  and  a28803a );
 a28813a <=( A234  and  A232 );
 a28814a <=( A203  and  a28813a );
 a28818a <=( A302  and  (not A299) );
 a28819a <=( A298  and  a28818a );
 a28820a <=( a28819a  and  a28814a );
 a28823a <=( (not A169)  and  (not A170) );
 a28827a <=( A200  and  (not A199) );
 a28828a <=( (not A168)  and  a28827a );
 a28829a <=( a28828a  and  a28823a );
 a28833a <=( A234  and  A232 );
 a28834a <=( A203  and  a28833a );
 a28838a <=( A302  and  A299 );
 a28839a <=( (not A298)  and  a28838a );
 a28840a <=( a28839a  and  a28834a );
 a28843a <=( (not A169)  and  (not A170) );
 a28847a <=( A200  and  (not A199) );
 a28848a <=( (not A168)  and  a28847a );
 a28849a <=( a28848a  and  a28843a );
 a28853a <=( A234  and  A232 );
 a28854a <=( A203  and  a28853a );
 a28858a <=( A269  and  A266 );
 a28859a <=( (not A265)  and  a28858a );
 a28860a <=( a28859a  and  a28854a );
 a28863a <=( (not A169)  and  (not A170) );
 a28867a <=( A200  and  (not A199) );
 a28868a <=( (not A168)  and  a28867a );
 a28869a <=( a28868a  and  a28863a );
 a28873a <=( A234  and  A232 );
 a28874a <=( A203  and  a28873a );
 a28878a <=( A269  and  (not A266) );
 a28879a <=( A265  and  a28878a );
 a28880a <=( a28879a  and  a28874a );
 a28883a <=( (not A169)  and  (not A170) );
 a28887a <=( A200  and  (not A199) );
 a28888a <=( (not A168)  and  a28887a );
 a28889a <=( a28888a  and  a28883a );
 a28893a <=( A234  and  A233 );
 a28894a <=( A203  and  a28893a );
 a28898a <=( A302  and  (not A299) );
 a28899a <=( A298  and  a28898a );
 a28900a <=( a28899a  and  a28894a );
 a28903a <=( (not A169)  and  (not A170) );
 a28907a <=( A200  and  (not A199) );
 a28908a <=( (not A168)  and  a28907a );
 a28909a <=( a28908a  and  a28903a );
 a28913a <=( A234  and  A233 );
 a28914a <=( A203  and  a28913a );
 a28918a <=( A302  and  A299 );
 a28919a <=( (not A298)  and  a28918a );
 a28920a <=( a28919a  and  a28914a );
 a28923a <=( (not A169)  and  (not A170) );
 a28927a <=( A200  and  (not A199) );
 a28928a <=( (not A168)  and  a28927a );
 a28929a <=( a28928a  and  a28923a );
 a28933a <=( A234  and  A233 );
 a28934a <=( A203  and  a28933a );
 a28938a <=( A269  and  A266 );
 a28939a <=( (not A265)  and  a28938a );
 a28940a <=( a28939a  and  a28934a );
 a28943a <=( (not A169)  and  (not A170) );
 a28947a <=( A200  and  (not A199) );
 a28948a <=( (not A168)  and  a28947a );
 a28949a <=( a28948a  and  a28943a );
 a28953a <=( A234  and  A233 );
 a28954a <=( A203  and  a28953a );
 a28958a <=( A269  and  (not A266) );
 a28959a <=( A265  and  a28958a );
 a28960a <=( a28959a  and  a28954a );
 a28963a <=( (not A169)  and  (not A170) );
 a28967a <=( A200  and  (not A199) );
 a28968a <=( (not A168)  and  a28967a );
 a28969a <=( a28968a  and  a28963a );
 a28973a <=( A233  and  (not A232) );
 a28974a <=( A203  and  a28973a );
 a28978a <=( A300  and  A299 );
 a28979a <=( A236  and  a28978a );
 a28980a <=( a28979a  and  a28974a );
 a28983a <=( (not A169)  and  (not A170) );
 a28987a <=( A200  and  (not A199) );
 a28988a <=( (not A168)  and  a28987a );
 a28989a <=( a28988a  and  a28983a );
 a28993a <=( A233  and  (not A232) );
 a28994a <=( A203  and  a28993a );
 a28998a <=( A300  and  A298 );
 a28999a <=( A236  and  a28998a );
 a29000a <=( a28999a  and  a28994a );
 a29003a <=( (not A169)  and  (not A170) );
 a29007a <=( A200  and  (not A199) );
 a29008a <=( (not A168)  and  a29007a );
 a29009a <=( a29008a  and  a29003a );
 a29013a <=( A233  and  (not A232) );
 a29014a <=( A203  and  a29013a );
 a29018a <=( A267  and  A265 );
 a29019a <=( A236  and  a29018a );
 a29020a <=( a29019a  and  a29014a );
 a29023a <=( (not A169)  and  (not A170) );
 a29027a <=( A200  and  (not A199) );
 a29028a <=( (not A168)  and  a29027a );
 a29029a <=( a29028a  and  a29023a );
 a29033a <=( A233  and  (not A232) );
 a29034a <=( A203  and  a29033a );
 a29038a <=( A267  and  A266 );
 a29039a <=( A236  and  a29038a );
 a29040a <=( a29039a  and  a29034a );
 a29043a <=( (not A169)  and  (not A170) );
 a29047a <=( A200  and  (not A199) );
 a29048a <=( (not A168)  and  a29047a );
 a29049a <=( a29048a  and  a29043a );
 a29053a <=( (not A233)  and  A232 );
 a29054a <=( A203  and  a29053a );
 a29058a <=( A300  and  A299 );
 a29059a <=( A236  and  a29058a );
 a29060a <=( a29059a  and  a29054a );
 a29063a <=( (not A169)  and  (not A170) );
 a29067a <=( A200  and  (not A199) );
 a29068a <=( (not A168)  and  a29067a );
 a29069a <=( a29068a  and  a29063a );
 a29073a <=( (not A233)  and  A232 );
 a29074a <=( A203  and  a29073a );
 a29078a <=( A300  and  A298 );
 a29079a <=( A236  and  a29078a );
 a29080a <=( a29079a  and  a29074a );
 a29083a <=( (not A169)  and  (not A170) );
 a29087a <=( A200  and  (not A199) );
 a29088a <=( (not A168)  and  a29087a );
 a29089a <=( a29088a  and  a29083a );
 a29093a <=( (not A233)  and  A232 );
 a29094a <=( A203  and  a29093a );
 a29098a <=( A267  and  A265 );
 a29099a <=( A236  and  a29098a );
 a29100a <=( a29099a  and  a29094a );
 a29103a <=( (not A169)  and  (not A170) );
 a29107a <=( A200  and  (not A199) );
 a29108a <=( (not A168)  and  a29107a );
 a29109a <=( a29108a  and  a29103a );
 a29113a <=( (not A233)  and  A232 );
 a29114a <=( A203  and  a29113a );
 a29118a <=( A267  and  A266 );
 a29119a <=( A236  and  a29118a );
 a29120a <=( a29119a  and  a29114a );
 a29123a <=( (not A169)  and  (not A170) );
 a29127a <=( (not A200)  and  A199 );
 a29128a <=( (not A168)  and  a29127a );
 a29129a <=( a29128a  and  a29123a );
 a29133a <=( A234  and  A232 );
 a29134a <=( A203  and  a29133a );
 a29138a <=( A302  and  (not A299) );
 a29139a <=( A298  and  a29138a );
 a29140a <=( a29139a  and  a29134a );
 a29143a <=( (not A169)  and  (not A170) );
 a29147a <=( (not A200)  and  A199 );
 a29148a <=( (not A168)  and  a29147a );
 a29149a <=( a29148a  and  a29143a );
 a29153a <=( A234  and  A232 );
 a29154a <=( A203  and  a29153a );
 a29158a <=( A302  and  A299 );
 a29159a <=( (not A298)  and  a29158a );
 a29160a <=( a29159a  and  a29154a );
 a29163a <=( (not A169)  and  (not A170) );
 a29167a <=( (not A200)  and  A199 );
 a29168a <=( (not A168)  and  a29167a );
 a29169a <=( a29168a  and  a29163a );
 a29173a <=( A234  and  A232 );
 a29174a <=( A203  and  a29173a );
 a29178a <=( A269  and  A266 );
 a29179a <=( (not A265)  and  a29178a );
 a29180a <=( a29179a  and  a29174a );
 a29183a <=( (not A169)  and  (not A170) );
 a29187a <=( (not A200)  and  A199 );
 a29188a <=( (not A168)  and  a29187a );
 a29189a <=( a29188a  and  a29183a );
 a29193a <=( A234  and  A232 );
 a29194a <=( A203  and  a29193a );
 a29198a <=( A269  and  (not A266) );
 a29199a <=( A265  and  a29198a );
 a29200a <=( a29199a  and  a29194a );
 a29203a <=( (not A169)  and  (not A170) );
 a29207a <=( (not A200)  and  A199 );
 a29208a <=( (not A168)  and  a29207a );
 a29209a <=( a29208a  and  a29203a );
 a29213a <=( A234  and  A233 );
 a29214a <=( A203  and  a29213a );
 a29218a <=( A302  and  (not A299) );
 a29219a <=( A298  and  a29218a );
 a29220a <=( a29219a  and  a29214a );
 a29223a <=( (not A169)  and  (not A170) );
 a29227a <=( (not A200)  and  A199 );
 a29228a <=( (not A168)  and  a29227a );
 a29229a <=( a29228a  and  a29223a );
 a29233a <=( A234  and  A233 );
 a29234a <=( A203  and  a29233a );
 a29238a <=( A302  and  A299 );
 a29239a <=( (not A298)  and  a29238a );
 a29240a <=( a29239a  and  a29234a );
 a29243a <=( (not A169)  and  (not A170) );
 a29247a <=( (not A200)  and  A199 );
 a29248a <=( (not A168)  and  a29247a );
 a29249a <=( a29248a  and  a29243a );
 a29253a <=( A234  and  A233 );
 a29254a <=( A203  and  a29253a );
 a29258a <=( A269  and  A266 );
 a29259a <=( (not A265)  and  a29258a );
 a29260a <=( a29259a  and  a29254a );
 a29263a <=( (not A169)  and  (not A170) );
 a29267a <=( (not A200)  and  A199 );
 a29268a <=( (not A168)  and  a29267a );
 a29269a <=( a29268a  and  a29263a );
 a29273a <=( A234  and  A233 );
 a29274a <=( A203  and  a29273a );
 a29278a <=( A269  and  (not A266) );
 a29279a <=( A265  and  a29278a );
 a29280a <=( a29279a  and  a29274a );
 a29283a <=( (not A169)  and  (not A170) );
 a29287a <=( (not A200)  and  A199 );
 a29288a <=( (not A168)  and  a29287a );
 a29289a <=( a29288a  and  a29283a );
 a29293a <=( A233  and  (not A232) );
 a29294a <=( A203  and  a29293a );
 a29298a <=( A300  and  A299 );
 a29299a <=( A236  and  a29298a );
 a29300a <=( a29299a  and  a29294a );
 a29303a <=( (not A169)  and  (not A170) );
 a29307a <=( (not A200)  and  A199 );
 a29308a <=( (not A168)  and  a29307a );
 a29309a <=( a29308a  and  a29303a );
 a29313a <=( A233  and  (not A232) );
 a29314a <=( A203  and  a29313a );
 a29318a <=( A300  and  A298 );
 a29319a <=( A236  and  a29318a );
 a29320a <=( a29319a  and  a29314a );
 a29323a <=( (not A169)  and  (not A170) );
 a29327a <=( (not A200)  and  A199 );
 a29328a <=( (not A168)  and  a29327a );
 a29329a <=( a29328a  and  a29323a );
 a29333a <=( A233  and  (not A232) );
 a29334a <=( A203  and  a29333a );
 a29338a <=( A267  and  A265 );
 a29339a <=( A236  and  a29338a );
 a29340a <=( a29339a  and  a29334a );
 a29343a <=( (not A169)  and  (not A170) );
 a29347a <=( (not A200)  and  A199 );
 a29348a <=( (not A168)  and  a29347a );
 a29349a <=( a29348a  and  a29343a );
 a29353a <=( A233  and  (not A232) );
 a29354a <=( A203  and  a29353a );
 a29358a <=( A267  and  A266 );
 a29359a <=( A236  and  a29358a );
 a29360a <=( a29359a  and  a29354a );
 a29363a <=( (not A169)  and  (not A170) );
 a29367a <=( (not A200)  and  A199 );
 a29368a <=( (not A168)  and  a29367a );
 a29369a <=( a29368a  and  a29363a );
 a29373a <=( (not A233)  and  A232 );
 a29374a <=( A203  and  a29373a );
 a29378a <=( A300  and  A299 );
 a29379a <=( A236  and  a29378a );
 a29380a <=( a29379a  and  a29374a );
 a29383a <=( (not A169)  and  (not A170) );
 a29387a <=( (not A200)  and  A199 );
 a29388a <=( (not A168)  and  a29387a );
 a29389a <=( a29388a  and  a29383a );
 a29393a <=( (not A233)  and  A232 );
 a29394a <=( A203  and  a29393a );
 a29398a <=( A300  and  A298 );
 a29399a <=( A236  and  a29398a );
 a29400a <=( a29399a  and  a29394a );
 a29403a <=( (not A169)  and  (not A170) );
 a29407a <=( (not A200)  and  A199 );
 a29408a <=( (not A168)  and  a29407a );
 a29409a <=( a29408a  and  a29403a );
 a29413a <=( (not A233)  and  A232 );
 a29414a <=( A203  and  a29413a );
 a29418a <=( A267  and  A265 );
 a29419a <=( A236  and  a29418a );
 a29420a <=( a29419a  and  a29414a );
 a29423a <=( (not A169)  and  (not A170) );
 a29427a <=( (not A200)  and  A199 );
 a29428a <=( (not A168)  and  a29427a );
 a29429a <=( a29428a  and  a29423a );
 a29433a <=( (not A233)  and  A232 );
 a29434a <=( A203  and  a29433a );
 a29438a <=( A267  and  A266 );
 a29439a <=( A236  and  a29438a );
 a29440a <=( a29439a  and  a29434a );
 a29444a <=( A199  and  A166 );
 a29445a <=( A168  and  a29444a );
 a29449a <=( (not A202)  and  (not A201) );
 a29450a <=( A200  and  a29449a );
 a29451a <=( a29450a  and  a29445a );
 a29455a <=( A236  and  A233 );
 a29456a <=( (not A232)  and  a29455a );
 a29460a <=( A302  and  (not A299) );
 a29461a <=( A298  and  a29460a );
 a29462a <=( a29461a  and  a29456a );
 a29466a <=( A199  and  A166 );
 a29467a <=( A168  and  a29466a );
 a29471a <=( (not A202)  and  (not A201) );
 a29472a <=( A200  and  a29471a );
 a29473a <=( a29472a  and  a29467a );
 a29477a <=( A236  and  A233 );
 a29478a <=( (not A232)  and  a29477a );
 a29482a <=( A302  and  A299 );
 a29483a <=( (not A298)  and  a29482a );
 a29484a <=( a29483a  and  a29478a );
 a29488a <=( A199  and  A166 );
 a29489a <=( A168  and  a29488a );
 a29493a <=( (not A202)  and  (not A201) );
 a29494a <=( A200  and  a29493a );
 a29495a <=( a29494a  and  a29489a );
 a29499a <=( A236  and  A233 );
 a29500a <=( (not A232)  and  a29499a );
 a29504a <=( A269  and  A266 );
 a29505a <=( (not A265)  and  a29504a );
 a29506a <=( a29505a  and  a29500a );
 a29510a <=( A199  and  A166 );
 a29511a <=( A168  and  a29510a );
 a29515a <=( (not A202)  and  (not A201) );
 a29516a <=( A200  and  a29515a );
 a29517a <=( a29516a  and  a29511a );
 a29521a <=( A236  and  A233 );
 a29522a <=( (not A232)  and  a29521a );
 a29526a <=( A269  and  (not A266) );
 a29527a <=( A265  and  a29526a );
 a29528a <=( a29527a  and  a29522a );
 a29532a <=( A199  and  A166 );
 a29533a <=( A168  and  a29532a );
 a29537a <=( (not A202)  and  (not A201) );
 a29538a <=( A200  and  a29537a );
 a29539a <=( a29538a  and  a29533a );
 a29543a <=( A236  and  (not A233) );
 a29544a <=( A232  and  a29543a );
 a29548a <=( A302  and  (not A299) );
 a29549a <=( A298  and  a29548a );
 a29550a <=( a29549a  and  a29544a );
 a29554a <=( A199  and  A166 );
 a29555a <=( A168  and  a29554a );
 a29559a <=( (not A202)  and  (not A201) );
 a29560a <=( A200  and  a29559a );
 a29561a <=( a29560a  and  a29555a );
 a29565a <=( A236  and  (not A233) );
 a29566a <=( A232  and  a29565a );
 a29570a <=( A302  and  A299 );
 a29571a <=( (not A298)  and  a29570a );
 a29572a <=( a29571a  and  a29566a );
 a29576a <=( A199  and  A166 );
 a29577a <=( A168  and  a29576a );
 a29581a <=( (not A202)  and  (not A201) );
 a29582a <=( A200  and  a29581a );
 a29583a <=( a29582a  and  a29577a );
 a29587a <=( A236  and  (not A233) );
 a29588a <=( A232  and  a29587a );
 a29592a <=( A269  and  A266 );
 a29593a <=( (not A265)  and  a29592a );
 a29594a <=( a29593a  and  a29588a );
 a29598a <=( A199  and  A166 );
 a29599a <=( A168  and  a29598a );
 a29603a <=( (not A202)  and  (not A201) );
 a29604a <=( A200  and  a29603a );
 a29605a <=( a29604a  and  a29599a );
 a29609a <=( A236  and  (not A233) );
 a29610a <=( A232  and  a29609a );
 a29614a <=( A269  and  (not A266) );
 a29615a <=( A265  and  a29614a );
 a29616a <=( a29615a  and  a29610a );
 a29620a <=( A199  and  A167 );
 a29621a <=( A168  and  a29620a );
 a29625a <=( (not A202)  and  (not A201) );
 a29626a <=( A200  and  a29625a );
 a29627a <=( a29626a  and  a29621a );
 a29631a <=( A236  and  A233 );
 a29632a <=( (not A232)  and  a29631a );
 a29636a <=( A302  and  (not A299) );
 a29637a <=( A298  and  a29636a );
 a29638a <=( a29637a  and  a29632a );
 a29642a <=( A199  and  A167 );
 a29643a <=( A168  and  a29642a );
 a29647a <=( (not A202)  and  (not A201) );
 a29648a <=( A200  and  a29647a );
 a29649a <=( a29648a  and  a29643a );
 a29653a <=( A236  and  A233 );
 a29654a <=( (not A232)  and  a29653a );
 a29658a <=( A302  and  A299 );
 a29659a <=( (not A298)  and  a29658a );
 a29660a <=( a29659a  and  a29654a );
 a29664a <=( A199  and  A167 );
 a29665a <=( A168  and  a29664a );
 a29669a <=( (not A202)  and  (not A201) );
 a29670a <=( A200  and  a29669a );
 a29671a <=( a29670a  and  a29665a );
 a29675a <=( A236  and  A233 );
 a29676a <=( (not A232)  and  a29675a );
 a29680a <=( A269  and  A266 );
 a29681a <=( (not A265)  and  a29680a );
 a29682a <=( a29681a  and  a29676a );
 a29686a <=( A199  and  A167 );
 a29687a <=( A168  and  a29686a );
 a29691a <=( (not A202)  and  (not A201) );
 a29692a <=( A200  and  a29691a );
 a29693a <=( a29692a  and  a29687a );
 a29697a <=( A236  and  A233 );
 a29698a <=( (not A232)  and  a29697a );
 a29702a <=( A269  and  (not A266) );
 a29703a <=( A265  and  a29702a );
 a29704a <=( a29703a  and  a29698a );
 a29708a <=( A199  and  A167 );
 a29709a <=( A168  and  a29708a );
 a29713a <=( (not A202)  and  (not A201) );
 a29714a <=( A200  and  a29713a );
 a29715a <=( a29714a  and  a29709a );
 a29719a <=( A236  and  (not A233) );
 a29720a <=( A232  and  a29719a );
 a29724a <=( A302  and  (not A299) );
 a29725a <=( A298  and  a29724a );
 a29726a <=( a29725a  and  a29720a );
 a29730a <=( A199  and  A167 );
 a29731a <=( A168  and  a29730a );
 a29735a <=( (not A202)  and  (not A201) );
 a29736a <=( A200  and  a29735a );
 a29737a <=( a29736a  and  a29731a );
 a29741a <=( A236  and  (not A233) );
 a29742a <=( A232  and  a29741a );
 a29746a <=( A302  and  A299 );
 a29747a <=( (not A298)  and  a29746a );
 a29748a <=( a29747a  and  a29742a );
 a29752a <=( A199  and  A167 );
 a29753a <=( A168  and  a29752a );
 a29757a <=( (not A202)  and  (not A201) );
 a29758a <=( A200  and  a29757a );
 a29759a <=( a29758a  and  a29753a );
 a29763a <=( A236  and  (not A233) );
 a29764a <=( A232  and  a29763a );
 a29768a <=( A269  and  A266 );
 a29769a <=( (not A265)  and  a29768a );
 a29770a <=( a29769a  and  a29764a );
 a29774a <=( A199  and  A167 );
 a29775a <=( A168  and  a29774a );
 a29779a <=( (not A202)  and  (not A201) );
 a29780a <=( A200  and  a29779a );
 a29781a <=( a29780a  and  a29775a );
 a29785a <=( A236  and  (not A233) );
 a29786a <=( A232  and  a29785a );
 a29790a <=( A269  and  (not A266) );
 a29791a <=( A265  and  a29790a );
 a29792a <=( a29791a  and  a29786a );
 a29796a <=( (not A166)  and  A167 );
 a29797a <=( A170  and  a29796a );
 a29801a <=( (not A203)  and  (not A202) );
 a29802a <=( (not A201)  and  a29801a );
 a29803a <=( a29802a  and  a29797a );
 a29807a <=( A236  and  A233 );
 a29808a <=( (not A232)  and  a29807a );
 a29812a <=( A302  and  (not A299) );
 a29813a <=( A298  and  a29812a );
 a29814a <=( a29813a  and  a29808a );
 a29818a <=( (not A166)  and  A167 );
 a29819a <=( A170  and  a29818a );
 a29823a <=( (not A203)  and  (not A202) );
 a29824a <=( (not A201)  and  a29823a );
 a29825a <=( a29824a  and  a29819a );
 a29829a <=( A236  and  A233 );
 a29830a <=( (not A232)  and  a29829a );
 a29834a <=( A302  and  A299 );
 a29835a <=( (not A298)  and  a29834a );
 a29836a <=( a29835a  and  a29830a );
 a29840a <=( (not A166)  and  A167 );
 a29841a <=( A170  and  a29840a );
 a29845a <=( (not A203)  and  (not A202) );
 a29846a <=( (not A201)  and  a29845a );
 a29847a <=( a29846a  and  a29841a );
 a29851a <=( A236  and  A233 );
 a29852a <=( (not A232)  and  a29851a );
 a29856a <=( A269  and  A266 );
 a29857a <=( (not A265)  and  a29856a );
 a29858a <=( a29857a  and  a29852a );
 a29862a <=( (not A166)  and  A167 );
 a29863a <=( A170  and  a29862a );
 a29867a <=( (not A203)  and  (not A202) );
 a29868a <=( (not A201)  and  a29867a );
 a29869a <=( a29868a  and  a29863a );
 a29873a <=( A236  and  A233 );
 a29874a <=( (not A232)  and  a29873a );
 a29878a <=( A269  and  (not A266) );
 a29879a <=( A265  and  a29878a );
 a29880a <=( a29879a  and  a29874a );
 a29884a <=( (not A166)  and  A167 );
 a29885a <=( A170  and  a29884a );
 a29889a <=( (not A203)  and  (not A202) );
 a29890a <=( (not A201)  and  a29889a );
 a29891a <=( a29890a  and  a29885a );
 a29895a <=( A236  and  (not A233) );
 a29896a <=( A232  and  a29895a );
 a29900a <=( A302  and  (not A299) );
 a29901a <=( A298  and  a29900a );
 a29902a <=( a29901a  and  a29896a );
 a29906a <=( (not A166)  and  A167 );
 a29907a <=( A170  and  a29906a );
 a29911a <=( (not A203)  and  (not A202) );
 a29912a <=( (not A201)  and  a29911a );
 a29913a <=( a29912a  and  a29907a );
 a29917a <=( A236  and  (not A233) );
 a29918a <=( A232  and  a29917a );
 a29922a <=( A302  and  A299 );
 a29923a <=( (not A298)  and  a29922a );
 a29924a <=( a29923a  and  a29918a );
 a29928a <=( (not A166)  and  A167 );
 a29929a <=( A170  and  a29928a );
 a29933a <=( (not A203)  and  (not A202) );
 a29934a <=( (not A201)  and  a29933a );
 a29935a <=( a29934a  and  a29929a );
 a29939a <=( A236  and  (not A233) );
 a29940a <=( A232  and  a29939a );
 a29944a <=( A269  and  A266 );
 a29945a <=( (not A265)  and  a29944a );
 a29946a <=( a29945a  and  a29940a );
 a29950a <=( (not A166)  and  A167 );
 a29951a <=( A170  and  a29950a );
 a29955a <=( (not A203)  and  (not A202) );
 a29956a <=( (not A201)  and  a29955a );
 a29957a <=( a29956a  and  a29951a );
 a29961a <=( A236  and  (not A233) );
 a29962a <=( A232  and  a29961a );
 a29966a <=( A269  and  (not A266) );
 a29967a <=( A265  and  a29966a );
 a29968a <=( a29967a  and  a29962a );
 a29972a <=( (not A166)  and  A167 );
 a29973a <=( A170  and  a29972a );
 a29977a <=( (not A201)  and  A200 );
 a29978a <=( A199  and  a29977a );
 a29979a <=( a29978a  and  a29973a );
 a29983a <=( A234  and  A232 );
 a29984a <=( (not A202)  and  a29983a );
 a29988a <=( A302  and  (not A299) );
 a29989a <=( A298  and  a29988a );
 a29990a <=( a29989a  and  a29984a );
 a29994a <=( (not A166)  and  A167 );
 a29995a <=( A170  and  a29994a );
 a29999a <=( (not A201)  and  A200 );
 a30000a <=( A199  and  a29999a );
 a30001a <=( a30000a  and  a29995a );
 a30005a <=( A234  and  A232 );
 a30006a <=( (not A202)  and  a30005a );
 a30010a <=( A302  and  A299 );
 a30011a <=( (not A298)  and  a30010a );
 a30012a <=( a30011a  and  a30006a );
 a30016a <=( (not A166)  and  A167 );
 a30017a <=( A170  and  a30016a );
 a30021a <=( (not A201)  and  A200 );
 a30022a <=( A199  and  a30021a );
 a30023a <=( a30022a  and  a30017a );
 a30027a <=( A234  and  A232 );
 a30028a <=( (not A202)  and  a30027a );
 a30032a <=( A269  and  A266 );
 a30033a <=( (not A265)  and  a30032a );
 a30034a <=( a30033a  and  a30028a );
 a30038a <=( (not A166)  and  A167 );
 a30039a <=( A170  and  a30038a );
 a30043a <=( (not A201)  and  A200 );
 a30044a <=( A199  and  a30043a );
 a30045a <=( a30044a  and  a30039a );
 a30049a <=( A234  and  A232 );
 a30050a <=( (not A202)  and  a30049a );
 a30054a <=( A269  and  (not A266) );
 a30055a <=( A265  and  a30054a );
 a30056a <=( a30055a  and  a30050a );
 a30060a <=( (not A166)  and  A167 );
 a30061a <=( A170  and  a30060a );
 a30065a <=( (not A201)  and  A200 );
 a30066a <=( A199  and  a30065a );
 a30067a <=( a30066a  and  a30061a );
 a30071a <=( A234  and  A233 );
 a30072a <=( (not A202)  and  a30071a );
 a30076a <=( A302  and  (not A299) );
 a30077a <=( A298  and  a30076a );
 a30078a <=( a30077a  and  a30072a );
 a30082a <=( (not A166)  and  A167 );
 a30083a <=( A170  and  a30082a );
 a30087a <=( (not A201)  and  A200 );
 a30088a <=( A199  and  a30087a );
 a30089a <=( a30088a  and  a30083a );
 a30093a <=( A234  and  A233 );
 a30094a <=( (not A202)  and  a30093a );
 a30098a <=( A302  and  A299 );
 a30099a <=( (not A298)  and  a30098a );
 a30100a <=( a30099a  and  a30094a );
 a30104a <=( (not A166)  and  A167 );
 a30105a <=( A170  and  a30104a );
 a30109a <=( (not A201)  and  A200 );
 a30110a <=( A199  and  a30109a );
 a30111a <=( a30110a  and  a30105a );
 a30115a <=( A234  and  A233 );
 a30116a <=( (not A202)  and  a30115a );
 a30120a <=( A269  and  A266 );
 a30121a <=( (not A265)  and  a30120a );
 a30122a <=( a30121a  and  a30116a );
 a30126a <=( (not A166)  and  A167 );
 a30127a <=( A170  and  a30126a );
 a30131a <=( (not A201)  and  A200 );
 a30132a <=( A199  and  a30131a );
 a30133a <=( a30132a  and  a30127a );
 a30137a <=( A234  and  A233 );
 a30138a <=( (not A202)  and  a30137a );
 a30142a <=( A269  and  (not A266) );
 a30143a <=( A265  and  a30142a );
 a30144a <=( a30143a  and  a30138a );
 a30148a <=( (not A166)  and  A167 );
 a30149a <=( A170  and  a30148a );
 a30153a <=( (not A201)  and  A200 );
 a30154a <=( A199  and  a30153a );
 a30155a <=( a30154a  and  a30149a );
 a30159a <=( A233  and  (not A232) );
 a30160a <=( (not A202)  and  a30159a );
 a30164a <=( A300  and  A299 );
 a30165a <=( A236  and  a30164a );
 a30166a <=( a30165a  and  a30160a );
 a30170a <=( (not A166)  and  A167 );
 a30171a <=( A170  and  a30170a );
 a30175a <=( (not A201)  and  A200 );
 a30176a <=( A199  and  a30175a );
 a30177a <=( a30176a  and  a30171a );
 a30181a <=( A233  and  (not A232) );
 a30182a <=( (not A202)  and  a30181a );
 a30186a <=( A300  and  A298 );
 a30187a <=( A236  and  a30186a );
 a30188a <=( a30187a  and  a30182a );
 a30192a <=( (not A166)  and  A167 );
 a30193a <=( A170  and  a30192a );
 a30197a <=( (not A201)  and  A200 );
 a30198a <=( A199  and  a30197a );
 a30199a <=( a30198a  and  a30193a );
 a30203a <=( A233  and  (not A232) );
 a30204a <=( (not A202)  and  a30203a );
 a30208a <=( A267  and  A265 );
 a30209a <=( A236  and  a30208a );
 a30210a <=( a30209a  and  a30204a );
 a30214a <=( (not A166)  and  A167 );
 a30215a <=( A170  and  a30214a );
 a30219a <=( (not A201)  and  A200 );
 a30220a <=( A199  and  a30219a );
 a30221a <=( a30220a  and  a30215a );
 a30225a <=( A233  and  (not A232) );
 a30226a <=( (not A202)  and  a30225a );
 a30230a <=( A267  and  A266 );
 a30231a <=( A236  and  a30230a );
 a30232a <=( a30231a  and  a30226a );
 a30236a <=( (not A166)  and  A167 );
 a30237a <=( A170  and  a30236a );
 a30241a <=( (not A201)  and  A200 );
 a30242a <=( A199  and  a30241a );
 a30243a <=( a30242a  and  a30237a );
 a30247a <=( (not A233)  and  A232 );
 a30248a <=( (not A202)  and  a30247a );
 a30252a <=( A300  and  A299 );
 a30253a <=( A236  and  a30252a );
 a30254a <=( a30253a  and  a30248a );
 a30258a <=( (not A166)  and  A167 );
 a30259a <=( A170  and  a30258a );
 a30263a <=( (not A201)  and  A200 );
 a30264a <=( A199  and  a30263a );
 a30265a <=( a30264a  and  a30259a );
 a30269a <=( (not A233)  and  A232 );
 a30270a <=( (not A202)  and  a30269a );
 a30274a <=( A300  and  A298 );
 a30275a <=( A236  and  a30274a );
 a30276a <=( a30275a  and  a30270a );
 a30280a <=( (not A166)  and  A167 );
 a30281a <=( A170  and  a30280a );
 a30285a <=( (not A201)  and  A200 );
 a30286a <=( A199  and  a30285a );
 a30287a <=( a30286a  and  a30281a );
 a30291a <=( (not A233)  and  A232 );
 a30292a <=( (not A202)  and  a30291a );
 a30296a <=( A267  and  A265 );
 a30297a <=( A236  and  a30296a );
 a30298a <=( a30297a  and  a30292a );
 a30302a <=( (not A166)  and  A167 );
 a30303a <=( A170  and  a30302a );
 a30307a <=( (not A201)  and  A200 );
 a30308a <=( A199  and  a30307a );
 a30309a <=( a30308a  and  a30303a );
 a30313a <=( (not A233)  and  A232 );
 a30314a <=( (not A202)  and  a30313a );
 a30318a <=( A267  and  A266 );
 a30319a <=( A236  and  a30318a );
 a30320a <=( a30319a  and  a30314a );
 a30324a <=( (not A166)  and  A167 );
 a30325a <=( A170  and  a30324a );
 a30329a <=( (not A202)  and  (not A200) );
 a30330a <=( (not A199)  and  a30329a );
 a30331a <=( a30330a  and  a30325a );
 a30335a <=( A236  and  A233 );
 a30336a <=( (not A232)  and  a30335a );
 a30340a <=( A302  and  (not A299) );
 a30341a <=( A298  and  a30340a );
 a30342a <=( a30341a  and  a30336a );
 a30346a <=( (not A166)  and  A167 );
 a30347a <=( A170  and  a30346a );
 a30351a <=( (not A202)  and  (not A200) );
 a30352a <=( (not A199)  and  a30351a );
 a30353a <=( a30352a  and  a30347a );
 a30357a <=( A236  and  A233 );
 a30358a <=( (not A232)  and  a30357a );
 a30362a <=( A302  and  A299 );
 a30363a <=( (not A298)  and  a30362a );
 a30364a <=( a30363a  and  a30358a );
 a30368a <=( (not A166)  and  A167 );
 a30369a <=( A170  and  a30368a );
 a30373a <=( (not A202)  and  (not A200) );
 a30374a <=( (not A199)  and  a30373a );
 a30375a <=( a30374a  and  a30369a );
 a30379a <=( A236  and  A233 );
 a30380a <=( (not A232)  and  a30379a );
 a30384a <=( A269  and  A266 );
 a30385a <=( (not A265)  and  a30384a );
 a30386a <=( a30385a  and  a30380a );
 a30390a <=( (not A166)  and  A167 );
 a30391a <=( A170  and  a30390a );
 a30395a <=( (not A202)  and  (not A200) );
 a30396a <=( (not A199)  and  a30395a );
 a30397a <=( a30396a  and  a30391a );
 a30401a <=( A236  and  A233 );
 a30402a <=( (not A232)  and  a30401a );
 a30406a <=( A269  and  (not A266) );
 a30407a <=( A265  and  a30406a );
 a30408a <=( a30407a  and  a30402a );
 a30412a <=( (not A166)  and  A167 );
 a30413a <=( A170  and  a30412a );
 a30417a <=( (not A202)  and  (not A200) );
 a30418a <=( (not A199)  and  a30417a );
 a30419a <=( a30418a  and  a30413a );
 a30423a <=( A236  and  (not A233) );
 a30424a <=( A232  and  a30423a );
 a30428a <=( A302  and  (not A299) );
 a30429a <=( A298  and  a30428a );
 a30430a <=( a30429a  and  a30424a );
 a30434a <=( (not A166)  and  A167 );
 a30435a <=( A170  and  a30434a );
 a30439a <=( (not A202)  and  (not A200) );
 a30440a <=( (not A199)  and  a30439a );
 a30441a <=( a30440a  and  a30435a );
 a30445a <=( A236  and  (not A233) );
 a30446a <=( A232  and  a30445a );
 a30450a <=( A302  and  A299 );
 a30451a <=( (not A298)  and  a30450a );
 a30452a <=( a30451a  and  a30446a );
 a30456a <=( (not A166)  and  A167 );
 a30457a <=( A170  and  a30456a );
 a30461a <=( (not A202)  and  (not A200) );
 a30462a <=( (not A199)  and  a30461a );
 a30463a <=( a30462a  and  a30457a );
 a30467a <=( A236  and  (not A233) );
 a30468a <=( A232  and  a30467a );
 a30472a <=( A269  and  A266 );
 a30473a <=( (not A265)  and  a30472a );
 a30474a <=( a30473a  and  a30468a );
 a30478a <=( (not A166)  and  A167 );
 a30479a <=( A170  and  a30478a );
 a30483a <=( (not A202)  and  (not A200) );
 a30484a <=( (not A199)  and  a30483a );
 a30485a <=( a30484a  and  a30479a );
 a30489a <=( A236  and  (not A233) );
 a30490a <=( A232  and  a30489a );
 a30494a <=( A269  and  (not A266) );
 a30495a <=( A265  and  a30494a );
 a30496a <=( a30495a  and  a30490a );
 a30500a <=( A166  and  (not A167) );
 a30501a <=( A170  and  a30500a );
 a30505a <=( (not A203)  and  (not A202) );
 a30506a <=( (not A201)  and  a30505a );
 a30507a <=( a30506a  and  a30501a );
 a30511a <=( A236  and  A233 );
 a30512a <=( (not A232)  and  a30511a );
 a30516a <=( A302  and  (not A299) );
 a30517a <=( A298  and  a30516a );
 a30518a <=( a30517a  and  a30512a );
 a30522a <=( A166  and  (not A167) );
 a30523a <=( A170  and  a30522a );
 a30527a <=( (not A203)  and  (not A202) );
 a30528a <=( (not A201)  and  a30527a );
 a30529a <=( a30528a  and  a30523a );
 a30533a <=( A236  and  A233 );
 a30534a <=( (not A232)  and  a30533a );
 a30538a <=( A302  and  A299 );
 a30539a <=( (not A298)  and  a30538a );
 a30540a <=( a30539a  and  a30534a );
 a30544a <=( A166  and  (not A167) );
 a30545a <=( A170  and  a30544a );
 a30549a <=( (not A203)  and  (not A202) );
 a30550a <=( (not A201)  and  a30549a );
 a30551a <=( a30550a  and  a30545a );
 a30555a <=( A236  and  A233 );
 a30556a <=( (not A232)  and  a30555a );
 a30560a <=( A269  and  A266 );
 a30561a <=( (not A265)  and  a30560a );
 a30562a <=( a30561a  and  a30556a );
 a30566a <=( A166  and  (not A167) );
 a30567a <=( A170  and  a30566a );
 a30571a <=( (not A203)  and  (not A202) );
 a30572a <=( (not A201)  and  a30571a );
 a30573a <=( a30572a  and  a30567a );
 a30577a <=( A236  and  A233 );
 a30578a <=( (not A232)  and  a30577a );
 a30582a <=( A269  and  (not A266) );
 a30583a <=( A265  and  a30582a );
 a30584a <=( a30583a  and  a30578a );
 a30588a <=( A166  and  (not A167) );
 a30589a <=( A170  and  a30588a );
 a30593a <=( (not A203)  and  (not A202) );
 a30594a <=( (not A201)  and  a30593a );
 a30595a <=( a30594a  and  a30589a );
 a30599a <=( A236  and  (not A233) );
 a30600a <=( A232  and  a30599a );
 a30604a <=( A302  and  (not A299) );
 a30605a <=( A298  and  a30604a );
 a30606a <=( a30605a  and  a30600a );
 a30610a <=( A166  and  (not A167) );
 a30611a <=( A170  and  a30610a );
 a30615a <=( (not A203)  and  (not A202) );
 a30616a <=( (not A201)  and  a30615a );
 a30617a <=( a30616a  and  a30611a );
 a30621a <=( A236  and  (not A233) );
 a30622a <=( A232  and  a30621a );
 a30626a <=( A302  and  A299 );
 a30627a <=( (not A298)  and  a30626a );
 a30628a <=( a30627a  and  a30622a );
 a30632a <=( A166  and  (not A167) );
 a30633a <=( A170  and  a30632a );
 a30637a <=( (not A203)  and  (not A202) );
 a30638a <=( (not A201)  and  a30637a );
 a30639a <=( a30638a  and  a30633a );
 a30643a <=( A236  and  (not A233) );
 a30644a <=( A232  and  a30643a );
 a30648a <=( A269  and  A266 );
 a30649a <=( (not A265)  and  a30648a );
 a30650a <=( a30649a  and  a30644a );
 a30654a <=( A166  and  (not A167) );
 a30655a <=( A170  and  a30654a );
 a30659a <=( (not A203)  and  (not A202) );
 a30660a <=( (not A201)  and  a30659a );
 a30661a <=( a30660a  and  a30655a );
 a30665a <=( A236  and  (not A233) );
 a30666a <=( A232  and  a30665a );
 a30670a <=( A269  and  (not A266) );
 a30671a <=( A265  and  a30670a );
 a30672a <=( a30671a  and  a30666a );
 a30676a <=( A166  and  (not A167) );
 a30677a <=( A170  and  a30676a );
 a30681a <=( (not A201)  and  A200 );
 a30682a <=( A199  and  a30681a );
 a30683a <=( a30682a  and  a30677a );
 a30687a <=( A234  and  A232 );
 a30688a <=( (not A202)  and  a30687a );
 a30692a <=( A302  and  (not A299) );
 a30693a <=( A298  and  a30692a );
 a30694a <=( a30693a  and  a30688a );
 a30698a <=( A166  and  (not A167) );
 a30699a <=( A170  and  a30698a );
 a30703a <=( (not A201)  and  A200 );
 a30704a <=( A199  and  a30703a );
 a30705a <=( a30704a  and  a30699a );
 a30709a <=( A234  and  A232 );
 a30710a <=( (not A202)  and  a30709a );
 a30714a <=( A302  and  A299 );
 a30715a <=( (not A298)  and  a30714a );
 a30716a <=( a30715a  and  a30710a );
 a30720a <=( A166  and  (not A167) );
 a30721a <=( A170  and  a30720a );
 a30725a <=( (not A201)  and  A200 );
 a30726a <=( A199  and  a30725a );
 a30727a <=( a30726a  and  a30721a );
 a30731a <=( A234  and  A232 );
 a30732a <=( (not A202)  and  a30731a );
 a30736a <=( A269  and  A266 );
 a30737a <=( (not A265)  and  a30736a );
 a30738a <=( a30737a  and  a30732a );
 a30742a <=( A166  and  (not A167) );
 a30743a <=( A170  and  a30742a );
 a30747a <=( (not A201)  and  A200 );
 a30748a <=( A199  and  a30747a );
 a30749a <=( a30748a  and  a30743a );
 a30753a <=( A234  and  A232 );
 a30754a <=( (not A202)  and  a30753a );
 a30758a <=( A269  and  (not A266) );
 a30759a <=( A265  and  a30758a );
 a30760a <=( a30759a  and  a30754a );
 a30764a <=( A166  and  (not A167) );
 a30765a <=( A170  and  a30764a );
 a30769a <=( (not A201)  and  A200 );
 a30770a <=( A199  and  a30769a );
 a30771a <=( a30770a  and  a30765a );
 a30775a <=( A234  and  A233 );
 a30776a <=( (not A202)  and  a30775a );
 a30780a <=( A302  and  (not A299) );
 a30781a <=( A298  and  a30780a );
 a30782a <=( a30781a  and  a30776a );
 a30786a <=( A166  and  (not A167) );
 a30787a <=( A170  and  a30786a );
 a30791a <=( (not A201)  and  A200 );
 a30792a <=( A199  and  a30791a );
 a30793a <=( a30792a  and  a30787a );
 a30797a <=( A234  and  A233 );
 a30798a <=( (not A202)  and  a30797a );
 a30802a <=( A302  and  A299 );
 a30803a <=( (not A298)  and  a30802a );
 a30804a <=( a30803a  and  a30798a );
 a30808a <=( A166  and  (not A167) );
 a30809a <=( A170  and  a30808a );
 a30813a <=( (not A201)  and  A200 );
 a30814a <=( A199  and  a30813a );
 a30815a <=( a30814a  and  a30809a );
 a30819a <=( A234  and  A233 );
 a30820a <=( (not A202)  and  a30819a );
 a30824a <=( A269  and  A266 );
 a30825a <=( (not A265)  and  a30824a );
 a30826a <=( a30825a  and  a30820a );
 a30830a <=( A166  and  (not A167) );
 a30831a <=( A170  and  a30830a );
 a30835a <=( (not A201)  and  A200 );
 a30836a <=( A199  and  a30835a );
 a30837a <=( a30836a  and  a30831a );
 a30841a <=( A234  and  A233 );
 a30842a <=( (not A202)  and  a30841a );
 a30846a <=( A269  and  (not A266) );
 a30847a <=( A265  and  a30846a );
 a30848a <=( a30847a  and  a30842a );
 a30852a <=( A166  and  (not A167) );
 a30853a <=( A170  and  a30852a );
 a30857a <=( (not A201)  and  A200 );
 a30858a <=( A199  and  a30857a );
 a30859a <=( a30858a  and  a30853a );
 a30863a <=( A233  and  (not A232) );
 a30864a <=( (not A202)  and  a30863a );
 a30868a <=( A300  and  A299 );
 a30869a <=( A236  and  a30868a );
 a30870a <=( a30869a  and  a30864a );
 a30874a <=( A166  and  (not A167) );
 a30875a <=( A170  and  a30874a );
 a30879a <=( (not A201)  and  A200 );
 a30880a <=( A199  and  a30879a );
 a30881a <=( a30880a  and  a30875a );
 a30885a <=( A233  and  (not A232) );
 a30886a <=( (not A202)  and  a30885a );
 a30890a <=( A300  and  A298 );
 a30891a <=( A236  and  a30890a );
 a30892a <=( a30891a  and  a30886a );
 a30896a <=( A166  and  (not A167) );
 a30897a <=( A170  and  a30896a );
 a30901a <=( (not A201)  and  A200 );
 a30902a <=( A199  and  a30901a );
 a30903a <=( a30902a  and  a30897a );
 a30907a <=( A233  and  (not A232) );
 a30908a <=( (not A202)  and  a30907a );
 a30912a <=( A267  and  A265 );
 a30913a <=( A236  and  a30912a );
 a30914a <=( a30913a  and  a30908a );
 a30918a <=( A166  and  (not A167) );
 a30919a <=( A170  and  a30918a );
 a30923a <=( (not A201)  and  A200 );
 a30924a <=( A199  and  a30923a );
 a30925a <=( a30924a  and  a30919a );
 a30929a <=( A233  and  (not A232) );
 a30930a <=( (not A202)  and  a30929a );
 a30934a <=( A267  and  A266 );
 a30935a <=( A236  and  a30934a );
 a30936a <=( a30935a  and  a30930a );
 a30940a <=( A166  and  (not A167) );
 a30941a <=( A170  and  a30940a );
 a30945a <=( (not A201)  and  A200 );
 a30946a <=( A199  and  a30945a );
 a30947a <=( a30946a  and  a30941a );
 a30951a <=( (not A233)  and  A232 );
 a30952a <=( (not A202)  and  a30951a );
 a30956a <=( A300  and  A299 );
 a30957a <=( A236  and  a30956a );
 a30958a <=( a30957a  and  a30952a );
 a30962a <=( A166  and  (not A167) );
 a30963a <=( A170  and  a30962a );
 a30967a <=( (not A201)  and  A200 );
 a30968a <=( A199  and  a30967a );
 a30969a <=( a30968a  and  a30963a );
 a30973a <=( (not A233)  and  A232 );
 a30974a <=( (not A202)  and  a30973a );
 a30978a <=( A300  and  A298 );
 a30979a <=( A236  and  a30978a );
 a30980a <=( a30979a  and  a30974a );
 a30984a <=( A166  and  (not A167) );
 a30985a <=( A170  and  a30984a );
 a30989a <=( (not A201)  and  A200 );
 a30990a <=( A199  and  a30989a );
 a30991a <=( a30990a  and  a30985a );
 a30995a <=( (not A233)  and  A232 );
 a30996a <=( (not A202)  and  a30995a );
 a31000a <=( A267  and  A265 );
 a31001a <=( A236  and  a31000a );
 a31002a <=( a31001a  and  a30996a );
 a31006a <=( A166  and  (not A167) );
 a31007a <=( A170  and  a31006a );
 a31011a <=( (not A201)  and  A200 );
 a31012a <=( A199  and  a31011a );
 a31013a <=( a31012a  and  a31007a );
 a31017a <=( (not A233)  and  A232 );
 a31018a <=( (not A202)  and  a31017a );
 a31022a <=( A267  and  A266 );
 a31023a <=( A236  and  a31022a );
 a31024a <=( a31023a  and  a31018a );
 a31028a <=( A166  and  (not A167) );
 a31029a <=( A170  and  a31028a );
 a31033a <=( (not A202)  and  (not A200) );
 a31034a <=( (not A199)  and  a31033a );
 a31035a <=( a31034a  and  a31029a );
 a31039a <=( A236  and  A233 );
 a31040a <=( (not A232)  and  a31039a );
 a31044a <=( A302  and  (not A299) );
 a31045a <=( A298  and  a31044a );
 a31046a <=( a31045a  and  a31040a );
 a31050a <=( A166  and  (not A167) );
 a31051a <=( A170  and  a31050a );
 a31055a <=( (not A202)  and  (not A200) );
 a31056a <=( (not A199)  and  a31055a );
 a31057a <=( a31056a  and  a31051a );
 a31061a <=( A236  and  A233 );
 a31062a <=( (not A232)  and  a31061a );
 a31066a <=( A302  and  A299 );
 a31067a <=( (not A298)  and  a31066a );
 a31068a <=( a31067a  and  a31062a );
 a31072a <=( A166  and  (not A167) );
 a31073a <=( A170  and  a31072a );
 a31077a <=( (not A202)  and  (not A200) );
 a31078a <=( (not A199)  and  a31077a );
 a31079a <=( a31078a  and  a31073a );
 a31083a <=( A236  and  A233 );
 a31084a <=( (not A232)  and  a31083a );
 a31088a <=( A269  and  A266 );
 a31089a <=( (not A265)  and  a31088a );
 a31090a <=( a31089a  and  a31084a );
 a31094a <=( A166  and  (not A167) );
 a31095a <=( A170  and  a31094a );
 a31099a <=( (not A202)  and  (not A200) );
 a31100a <=( (not A199)  and  a31099a );
 a31101a <=( a31100a  and  a31095a );
 a31105a <=( A236  and  A233 );
 a31106a <=( (not A232)  and  a31105a );
 a31110a <=( A269  and  (not A266) );
 a31111a <=( A265  and  a31110a );
 a31112a <=( a31111a  and  a31106a );
 a31116a <=( A166  and  (not A167) );
 a31117a <=( A170  and  a31116a );
 a31121a <=( (not A202)  and  (not A200) );
 a31122a <=( (not A199)  and  a31121a );
 a31123a <=( a31122a  and  a31117a );
 a31127a <=( A236  and  (not A233) );
 a31128a <=( A232  and  a31127a );
 a31132a <=( A302  and  (not A299) );
 a31133a <=( A298  and  a31132a );
 a31134a <=( a31133a  and  a31128a );
 a31138a <=( A166  and  (not A167) );
 a31139a <=( A170  and  a31138a );
 a31143a <=( (not A202)  and  (not A200) );
 a31144a <=( (not A199)  and  a31143a );
 a31145a <=( a31144a  and  a31139a );
 a31149a <=( A236  and  (not A233) );
 a31150a <=( A232  and  a31149a );
 a31154a <=( A302  and  A299 );
 a31155a <=( (not A298)  and  a31154a );
 a31156a <=( a31155a  and  a31150a );
 a31160a <=( A166  and  (not A167) );
 a31161a <=( A170  and  a31160a );
 a31165a <=( (not A202)  and  (not A200) );
 a31166a <=( (not A199)  and  a31165a );
 a31167a <=( a31166a  and  a31161a );
 a31171a <=( A236  and  (not A233) );
 a31172a <=( A232  and  a31171a );
 a31176a <=( A269  and  A266 );
 a31177a <=( (not A265)  and  a31176a );
 a31178a <=( a31177a  and  a31172a );
 a31182a <=( A166  and  (not A167) );
 a31183a <=( A170  and  a31182a );
 a31187a <=( (not A202)  and  (not A200) );
 a31188a <=( (not A199)  and  a31187a );
 a31189a <=( a31188a  and  a31183a );
 a31193a <=( A236  and  (not A233) );
 a31194a <=( A232  and  a31193a );
 a31198a <=( A269  and  (not A266) );
 a31199a <=( A265  and  a31198a );
 a31200a <=( a31199a  and  a31194a );
 a31204a <=( (not A166)  and  (not A167) );
 a31205a <=( (not A169)  and  a31204a );
 a31209a <=( A203  and  A200 );
 a31210a <=( (not A199)  and  a31209a );
 a31211a <=( a31210a  and  a31205a );
 a31215a <=( A236  and  A233 );
 a31216a <=( (not A232)  and  a31215a );
 a31220a <=( A302  and  (not A299) );
 a31221a <=( A298  and  a31220a );
 a31222a <=( a31221a  and  a31216a );
 a31226a <=( (not A166)  and  (not A167) );
 a31227a <=( (not A169)  and  a31226a );
 a31231a <=( A203  and  A200 );
 a31232a <=( (not A199)  and  a31231a );
 a31233a <=( a31232a  and  a31227a );
 a31237a <=( A236  and  A233 );
 a31238a <=( (not A232)  and  a31237a );
 a31242a <=( A302  and  A299 );
 a31243a <=( (not A298)  and  a31242a );
 a31244a <=( a31243a  and  a31238a );
 a31248a <=( (not A166)  and  (not A167) );
 a31249a <=( (not A169)  and  a31248a );
 a31253a <=( A203  and  A200 );
 a31254a <=( (not A199)  and  a31253a );
 a31255a <=( a31254a  and  a31249a );
 a31259a <=( A236  and  A233 );
 a31260a <=( (not A232)  and  a31259a );
 a31264a <=( A269  and  A266 );
 a31265a <=( (not A265)  and  a31264a );
 a31266a <=( a31265a  and  a31260a );
 a31270a <=( (not A166)  and  (not A167) );
 a31271a <=( (not A169)  and  a31270a );
 a31275a <=( A203  and  A200 );
 a31276a <=( (not A199)  and  a31275a );
 a31277a <=( a31276a  and  a31271a );
 a31281a <=( A236  and  A233 );
 a31282a <=( (not A232)  and  a31281a );
 a31286a <=( A269  and  (not A266) );
 a31287a <=( A265  and  a31286a );
 a31288a <=( a31287a  and  a31282a );
 a31292a <=( (not A166)  and  (not A167) );
 a31293a <=( (not A169)  and  a31292a );
 a31297a <=( A203  and  A200 );
 a31298a <=( (not A199)  and  a31297a );
 a31299a <=( a31298a  and  a31293a );
 a31303a <=( A236  and  (not A233) );
 a31304a <=( A232  and  a31303a );
 a31308a <=( A302  and  (not A299) );
 a31309a <=( A298  and  a31308a );
 a31310a <=( a31309a  and  a31304a );
 a31314a <=( (not A166)  and  (not A167) );
 a31315a <=( (not A169)  and  a31314a );
 a31319a <=( A203  and  A200 );
 a31320a <=( (not A199)  and  a31319a );
 a31321a <=( a31320a  and  a31315a );
 a31325a <=( A236  and  (not A233) );
 a31326a <=( A232  and  a31325a );
 a31330a <=( A302  and  A299 );
 a31331a <=( (not A298)  and  a31330a );
 a31332a <=( a31331a  and  a31326a );
 a31336a <=( (not A166)  and  (not A167) );
 a31337a <=( (not A169)  and  a31336a );
 a31341a <=( A203  and  A200 );
 a31342a <=( (not A199)  and  a31341a );
 a31343a <=( a31342a  and  a31337a );
 a31347a <=( A236  and  (not A233) );
 a31348a <=( A232  and  a31347a );
 a31352a <=( A269  and  A266 );
 a31353a <=( (not A265)  and  a31352a );
 a31354a <=( a31353a  and  a31348a );
 a31358a <=( (not A166)  and  (not A167) );
 a31359a <=( (not A169)  and  a31358a );
 a31363a <=( A203  and  A200 );
 a31364a <=( (not A199)  and  a31363a );
 a31365a <=( a31364a  and  a31359a );
 a31369a <=( A236  and  (not A233) );
 a31370a <=( A232  and  a31369a );
 a31374a <=( A269  and  (not A266) );
 a31375a <=( A265  and  a31374a );
 a31376a <=( a31375a  and  a31370a );
 a31380a <=( (not A166)  and  (not A167) );
 a31381a <=( (not A169)  and  a31380a );
 a31385a <=( A203  and  (not A200) );
 a31386a <=( A199  and  a31385a );
 a31387a <=( a31386a  and  a31381a );
 a31391a <=( A236  and  A233 );
 a31392a <=( (not A232)  and  a31391a );
 a31396a <=( A302  and  (not A299) );
 a31397a <=( A298  and  a31396a );
 a31398a <=( a31397a  and  a31392a );
 a31402a <=( (not A166)  and  (not A167) );
 a31403a <=( (not A169)  and  a31402a );
 a31407a <=( A203  and  (not A200) );
 a31408a <=( A199  and  a31407a );
 a31409a <=( a31408a  and  a31403a );
 a31413a <=( A236  and  A233 );
 a31414a <=( (not A232)  and  a31413a );
 a31418a <=( A302  and  A299 );
 a31419a <=( (not A298)  and  a31418a );
 a31420a <=( a31419a  and  a31414a );
 a31424a <=( (not A166)  and  (not A167) );
 a31425a <=( (not A169)  and  a31424a );
 a31429a <=( A203  and  (not A200) );
 a31430a <=( A199  and  a31429a );
 a31431a <=( a31430a  and  a31425a );
 a31435a <=( A236  and  A233 );
 a31436a <=( (not A232)  and  a31435a );
 a31440a <=( A269  and  A266 );
 a31441a <=( (not A265)  and  a31440a );
 a31442a <=( a31441a  and  a31436a );
 a31446a <=( (not A166)  and  (not A167) );
 a31447a <=( (not A169)  and  a31446a );
 a31451a <=( A203  and  (not A200) );
 a31452a <=( A199  and  a31451a );
 a31453a <=( a31452a  and  a31447a );
 a31457a <=( A236  and  A233 );
 a31458a <=( (not A232)  and  a31457a );
 a31462a <=( A269  and  (not A266) );
 a31463a <=( A265  and  a31462a );
 a31464a <=( a31463a  and  a31458a );
 a31468a <=( (not A166)  and  (not A167) );
 a31469a <=( (not A169)  and  a31468a );
 a31473a <=( A203  and  (not A200) );
 a31474a <=( A199  and  a31473a );
 a31475a <=( a31474a  and  a31469a );
 a31479a <=( A236  and  (not A233) );
 a31480a <=( A232  and  a31479a );
 a31484a <=( A302  and  (not A299) );
 a31485a <=( A298  and  a31484a );
 a31486a <=( a31485a  and  a31480a );
 a31490a <=( (not A166)  and  (not A167) );
 a31491a <=( (not A169)  and  a31490a );
 a31495a <=( A203  and  (not A200) );
 a31496a <=( A199  and  a31495a );
 a31497a <=( a31496a  and  a31491a );
 a31501a <=( A236  and  (not A233) );
 a31502a <=( A232  and  a31501a );
 a31506a <=( A302  and  A299 );
 a31507a <=( (not A298)  and  a31506a );
 a31508a <=( a31507a  and  a31502a );
 a31512a <=( (not A166)  and  (not A167) );
 a31513a <=( (not A169)  and  a31512a );
 a31517a <=( A203  and  (not A200) );
 a31518a <=( A199  and  a31517a );
 a31519a <=( a31518a  and  a31513a );
 a31523a <=( A236  and  (not A233) );
 a31524a <=( A232  and  a31523a );
 a31528a <=( A269  and  A266 );
 a31529a <=( (not A265)  and  a31528a );
 a31530a <=( a31529a  and  a31524a );
 a31534a <=( (not A166)  and  (not A167) );
 a31535a <=( (not A169)  and  a31534a );
 a31539a <=( A203  and  (not A200) );
 a31540a <=( A199  and  a31539a );
 a31541a <=( a31540a  and  a31535a );
 a31545a <=( A236  and  (not A233) );
 a31546a <=( A232  and  a31545a );
 a31550a <=( A269  and  (not A266) );
 a31551a <=( A265  and  a31550a );
 a31552a <=( a31551a  and  a31546a );
 a31556a <=( A167  and  (not A168) );
 a31557a <=( (not A169)  and  a31556a );
 a31561a <=( A201  and  A199 );
 a31562a <=( A166  and  a31561a );
 a31563a <=( a31562a  and  a31557a );
 a31567a <=( A236  and  A233 );
 a31568a <=( (not A232)  and  a31567a );
 a31572a <=( A302  and  (not A299) );
 a31573a <=( A298  and  a31572a );
 a31574a <=( a31573a  and  a31568a );
 a31578a <=( A167  and  (not A168) );
 a31579a <=( (not A169)  and  a31578a );
 a31583a <=( A201  and  A199 );
 a31584a <=( A166  and  a31583a );
 a31585a <=( a31584a  and  a31579a );
 a31589a <=( A236  and  A233 );
 a31590a <=( (not A232)  and  a31589a );
 a31594a <=( A302  and  A299 );
 a31595a <=( (not A298)  and  a31594a );
 a31596a <=( a31595a  and  a31590a );
 a31600a <=( A167  and  (not A168) );
 a31601a <=( (not A169)  and  a31600a );
 a31605a <=( A201  and  A199 );
 a31606a <=( A166  and  a31605a );
 a31607a <=( a31606a  and  a31601a );
 a31611a <=( A236  and  A233 );
 a31612a <=( (not A232)  and  a31611a );
 a31616a <=( A269  and  A266 );
 a31617a <=( (not A265)  and  a31616a );
 a31618a <=( a31617a  and  a31612a );
 a31622a <=( A167  and  (not A168) );
 a31623a <=( (not A169)  and  a31622a );
 a31627a <=( A201  and  A199 );
 a31628a <=( A166  and  a31627a );
 a31629a <=( a31628a  and  a31623a );
 a31633a <=( A236  and  A233 );
 a31634a <=( (not A232)  and  a31633a );
 a31638a <=( A269  and  (not A266) );
 a31639a <=( A265  and  a31638a );
 a31640a <=( a31639a  and  a31634a );
 a31644a <=( A167  and  (not A168) );
 a31645a <=( (not A169)  and  a31644a );
 a31649a <=( A201  and  A199 );
 a31650a <=( A166  and  a31649a );
 a31651a <=( a31650a  and  a31645a );
 a31655a <=( A236  and  (not A233) );
 a31656a <=( A232  and  a31655a );
 a31660a <=( A302  and  (not A299) );
 a31661a <=( A298  and  a31660a );
 a31662a <=( a31661a  and  a31656a );
 a31666a <=( A167  and  (not A168) );
 a31667a <=( (not A169)  and  a31666a );
 a31671a <=( A201  and  A199 );
 a31672a <=( A166  and  a31671a );
 a31673a <=( a31672a  and  a31667a );
 a31677a <=( A236  and  (not A233) );
 a31678a <=( A232  and  a31677a );
 a31682a <=( A302  and  A299 );
 a31683a <=( (not A298)  and  a31682a );
 a31684a <=( a31683a  and  a31678a );
 a31688a <=( A167  and  (not A168) );
 a31689a <=( (not A169)  and  a31688a );
 a31693a <=( A201  and  A199 );
 a31694a <=( A166  and  a31693a );
 a31695a <=( a31694a  and  a31689a );
 a31699a <=( A236  and  (not A233) );
 a31700a <=( A232  and  a31699a );
 a31704a <=( A269  and  A266 );
 a31705a <=( (not A265)  and  a31704a );
 a31706a <=( a31705a  and  a31700a );
 a31710a <=( A167  and  (not A168) );
 a31711a <=( (not A169)  and  a31710a );
 a31715a <=( A201  and  A199 );
 a31716a <=( A166  and  a31715a );
 a31717a <=( a31716a  and  a31711a );
 a31721a <=( A236  and  (not A233) );
 a31722a <=( A232  and  a31721a );
 a31726a <=( A269  and  (not A266) );
 a31727a <=( A265  and  a31726a );
 a31728a <=( a31727a  and  a31722a );
 a31732a <=( A167  and  (not A168) );
 a31733a <=( (not A169)  and  a31732a );
 a31737a <=( A201  and  A200 );
 a31738a <=( A166  and  a31737a );
 a31739a <=( a31738a  and  a31733a );
 a31743a <=( A236  and  A233 );
 a31744a <=( (not A232)  and  a31743a );
 a31748a <=( A302  and  (not A299) );
 a31749a <=( A298  and  a31748a );
 a31750a <=( a31749a  and  a31744a );
 a31754a <=( A167  and  (not A168) );
 a31755a <=( (not A169)  and  a31754a );
 a31759a <=( A201  and  A200 );
 a31760a <=( A166  and  a31759a );
 a31761a <=( a31760a  and  a31755a );
 a31765a <=( A236  and  A233 );
 a31766a <=( (not A232)  and  a31765a );
 a31770a <=( A302  and  A299 );
 a31771a <=( (not A298)  and  a31770a );
 a31772a <=( a31771a  and  a31766a );
 a31776a <=( A167  and  (not A168) );
 a31777a <=( (not A169)  and  a31776a );
 a31781a <=( A201  and  A200 );
 a31782a <=( A166  and  a31781a );
 a31783a <=( a31782a  and  a31777a );
 a31787a <=( A236  and  A233 );
 a31788a <=( (not A232)  and  a31787a );
 a31792a <=( A269  and  A266 );
 a31793a <=( (not A265)  and  a31792a );
 a31794a <=( a31793a  and  a31788a );
 a31798a <=( A167  and  (not A168) );
 a31799a <=( (not A169)  and  a31798a );
 a31803a <=( A201  and  A200 );
 a31804a <=( A166  and  a31803a );
 a31805a <=( a31804a  and  a31799a );
 a31809a <=( A236  and  A233 );
 a31810a <=( (not A232)  and  a31809a );
 a31814a <=( A269  and  (not A266) );
 a31815a <=( A265  and  a31814a );
 a31816a <=( a31815a  and  a31810a );
 a31820a <=( A167  and  (not A168) );
 a31821a <=( (not A169)  and  a31820a );
 a31825a <=( A201  and  A200 );
 a31826a <=( A166  and  a31825a );
 a31827a <=( a31826a  and  a31821a );
 a31831a <=( A236  and  (not A233) );
 a31832a <=( A232  and  a31831a );
 a31836a <=( A302  and  (not A299) );
 a31837a <=( A298  and  a31836a );
 a31838a <=( a31837a  and  a31832a );
 a31842a <=( A167  and  (not A168) );
 a31843a <=( (not A169)  and  a31842a );
 a31847a <=( A201  and  A200 );
 a31848a <=( A166  and  a31847a );
 a31849a <=( a31848a  and  a31843a );
 a31853a <=( A236  and  (not A233) );
 a31854a <=( A232  and  a31853a );
 a31858a <=( A302  and  A299 );
 a31859a <=( (not A298)  and  a31858a );
 a31860a <=( a31859a  and  a31854a );
 a31864a <=( A167  and  (not A168) );
 a31865a <=( (not A169)  and  a31864a );
 a31869a <=( A201  and  A200 );
 a31870a <=( A166  and  a31869a );
 a31871a <=( a31870a  and  a31865a );
 a31875a <=( A236  and  (not A233) );
 a31876a <=( A232  and  a31875a );
 a31880a <=( A269  and  A266 );
 a31881a <=( (not A265)  and  a31880a );
 a31882a <=( a31881a  and  a31876a );
 a31886a <=( A167  and  (not A168) );
 a31887a <=( (not A169)  and  a31886a );
 a31891a <=( A201  and  A200 );
 a31892a <=( A166  and  a31891a );
 a31893a <=( a31892a  and  a31887a );
 a31897a <=( A236  and  (not A233) );
 a31898a <=( A232  and  a31897a );
 a31902a <=( A269  and  (not A266) );
 a31903a <=( A265  and  a31902a );
 a31904a <=( a31903a  and  a31898a );
 a31908a <=( A167  and  (not A168) );
 a31909a <=( (not A169)  and  a31908a );
 a31913a <=( A200  and  (not A199) );
 a31914a <=( A166  and  a31913a );
 a31915a <=( a31914a  and  a31909a );
 a31919a <=( A234  and  A232 );
 a31920a <=( A203  and  a31919a );
 a31924a <=( A302  and  (not A299) );
 a31925a <=( A298  and  a31924a );
 a31926a <=( a31925a  and  a31920a );
 a31930a <=( A167  and  (not A168) );
 a31931a <=( (not A169)  and  a31930a );
 a31935a <=( A200  and  (not A199) );
 a31936a <=( A166  and  a31935a );
 a31937a <=( a31936a  and  a31931a );
 a31941a <=( A234  and  A232 );
 a31942a <=( A203  and  a31941a );
 a31946a <=( A302  and  A299 );
 a31947a <=( (not A298)  and  a31946a );
 a31948a <=( a31947a  and  a31942a );
 a31952a <=( A167  and  (not A168) );
 a31953a <=( (not A169)  and  a31952a );
 a31957a <=( A200  and  (not A199) );
 a31958a <=( A166  and  a31957a );
 a31959a <=( a31958a  and  a31953a );
 a31963a <=( A234  and  A232 );
 a31964a <=( A203  and  a31963a );
 a31968a <=( A269  and  A266 );
 a31969a <=( (not A265)  and  a31968a );
 a31970a <=( a31969a  and  a31964a );
 a31974a <=( A167  and  (not A168) );
 a31975a <=( (not A169)  and  a31974a );
 a31979a <=( A200  and  (not A199) );
 a31980a <=( A166  and  a31979a );
 a31981a <=( a31980a  and  a31975a );
 a31985a <=( A234  and  A232 );
 a31986a <=( A203  and  a31985a );
 a31990a <=( A269  and  (not A266) );
 a31991a <=( A265  and  a31990a );
 a31992a <=( a31991a  and  a31986a );
 a31996a <=( A167  and  (not A168) );
 a31997a <=( (not A169)  and  a31996a );
 a32001a <=( A200  and  (not A199) );
 a32002a <=( A166  and  a32001a );
 a32003a <=( a32002a  and  a31997a );
 a32007a <=( A234  and  A233 );
 a32008a <=( A203  and  a32007a );
 a32012a <=( A302  and  (not A299) );
 a32013a <=( A298  and  a32012a );
 a32014a <=( a32013a  and  a32008a );
 a32018a <=( A167  and  (not A168) );
 a32019a <=( (not A169)  and  a32018a );
 a32023a <=( A200  and  (not A199) );
 a32024a <=( A166  and  a32023a );
 a32025a <=( a32024a  and  a32019a );
 a32029a <=( A234  and  A233 );
 a32030a <=( A203  and  a32029a );
 a32034a <=( A302  and  A299 );
 a32035a <=( (not A298)  and  a32034a );
 a32036a <=( a32035a  and  a32030a );
 a32040a <=( A167  and  (not A168) );
 a32041a <=( (not A169)  and  a32040a );
 a32045a <=( A200  and  (not A199) );
 a32046a <=( A166  and  a32045a );
 a32047a <=( a32046a  and  a32041a );
 a32051a <=( A234  and  A233 );
 a32052a <=( A203  and  a32051a );
 a32056a <=( A269  and  A266 );
 a32057a <=( (not A265)  and  a32056a );
 a32058a <=( a32057a  and  a32052a );
 a32062a <=( A167  and  (not A168) );
 a32063a <=( (not A169)  and  a32062a );
 a32067a <=( A200  and  (not A199) );
 a32068a <=( A166  and  a32067a );
 a32069a <=( a32068a  and  a32063a );
 a32073a <=( A234  and  A233 );
 a32074a <=( A203  and  a32073a );
 a32078a <=( A269  and  (not A266) );
 a32079a <=( A265  and  a32078a );
 a32080a <=( a32079a  and  a32074a );
 a32084a <=( A167  and  (not A168) );
 a32085a <=( (not A169)  and  a32084a );
 a32089a <=( A200  and  (not A199) );
 a32090a <=( A166  and  a32089a );
 a32091a <=( a32090a  and  a32085a );
 a32095a <=( A233  and  (not A232) );
 a32096a <=( A203  and  a32095a );
 a32100a <=( A300  and  A299 );
 a32101a <=( A236  and  a32100a );
 a32102a <=( a32101a  and  a32096a );
 a32106a <=( A167  and  (not A168) );
 a32107a <=( (not A169)  and  a32106a );
 a32111a <=( A200  and  (not A199) );
 a32112a <=( A166  and  a32111a );
 a32113a <=( a32112a  and  a32107a );
 a32117a <=( A233  and  (not A232) );
 a32118a <=( A203  and  a32117a );
 a32122a <=( A300  and  A298 );
 a32123a <=( A236  and  a32122a );
 a32124a <=( a32123a  and  a32118a );
 a32128a <=( A167  and  (not A168) );
 a32129a <=( (not A169)  and  a32128a );
 a32133a <=( A200  and  (not A199) );
 a32134a <=( A166  and  a32133a );
 a32135a <=( a32134a  and  a32129a );
 a32139a <=( A233  and  (not A232) );
 a32140a <=( A203  and  a32139a );
 a32144a <=( A267  and  A265 );
 a32145a <=( A236  and  a32144a );
 a32146a <=( a32145a  and  a32140a );
 a32150a <=( A167  and  (not A168) );
 a32151a <=( (not A169)  and  a32150a );
 a32155a <=( A200  and  (not A199) );
 a32156a <=( A166  and  a32155a );
 a32157a <=( a32156a  and  a32151a );
 a32161a <=( A233  and  (not A232) );
 a32162a <=( A203  and  a32161a );
 a32166a <=( A267  and  A266 );
 a32167a <=( A236  and  a32166a );
 a32168a <=( a32167a  and  a32162a );
 a32172a <=( A167  and  (not A168) );
 a32173a <=( (not A169)  and  a32172a );
 a32177a <=( A200  and  (not A199) );
 a32178a <=( A166  and  a32177a );
 a32179a <=( a32178a  and  a32173a );
 a32183a <=( (not A233)  and  A232 );
 a32184a <=( A203  and  a32183a );
 a32188a <=( A300  and  A299 );
 a32189a <=( A236  and  a32188a );
 a32190a <=( a32189a  and  a32184a );
 a32194a <=( A167  and  (not A168) );
 a32195a <=( (not A169)  and  a32194a );
 a32199a <=( A200  and  (not A199) );
 a32200a <=( A166  and  a32199a );
 a32201a <=( a32200a  and  a32195a );
 a32205a <=( (not A233)  and  A232 );
 a32206a <=( A203  and  a32205a );
 a32210a <=( A300  and  A298 );
 a32211a <=( A236  and  a32210a );
 a32212a <=( a32211a  and  a32206a );
 a32216a <=( A167  and  (not A168) );
 a32217a <=( (not A169)  and  a32216a );
 a32221a <=( A200  and  (not A199) );
 a32222a <=( A166  and  a32221a );
 a32223a <=( a32222a  and  a32217a );
 a32227a <=( (not A233)  and  A232 );
 a32228a <=( A203  and  a32227a );
 a32232a <=( A267  and  A265 );
 a32233a <=( A236  and  a32232a );
 a32234a <=( a32233a  and  a32228a );
 a32238a <=( A167  and  (not A168) );
 a32239a <=( (not A169)  and  a32238a );
 a32243a <=( A200  and  (not A199) );
 a32244a <=( A166  and  a32243a );
 a32245a <=( a32244a  and  a32239a );
 a32249a <=( (not A233)  and  A232 );
 a32250a <=( A203  and  a32249a );
 a32254a <=( A267  and  A266 );
 a32255a <=( A236  and  a32254a );
 a32256a <=( a32255a  and  a32250a );
 a32260a <=( A167  and  (not A168) );
 a32261a <=( (not A169)  and  a32260a );
 a32265a <=( (not A200)  and  A199 );
 a32266a <=( A166  and  a32265a );
 a32267a <=( a32266a  and  a32261a );
 a32271a <=( A234  and  A232 );
 a32272a <=( A203  and  a32271a );
 a32276a <=( A302  and  (not A299) );
 a32277a <=( A298  and  a32276a );
 a32278a <=( a32277a  and  a32272a );
 a32282a <=( A167  and  (not A168) );
 a32283a <=( (not A169)  and  a32282a );
 a32287a <=( (not A200)  and  A199 );
 a32288a <=( A166  and  a32287a );
 a32289a <=( a32288a  and  a32283a );
 a32293a <=( A234  and  A232 );
 a32294a <=( A203  and  a32293a );
 a32298a <=( A302  and  A299 );
 a32299a <=( (not A298)  and  a32298a );
 a32300a <=( a32299a  and  a32294a );
 a32304a <=( A167  and  (not A168) );
 a32305a <=( (not A169)  and  a32304a );
 a32309a <=( (not A200)  and  A199 );
 a32310a <=( A166  and  a32309a );
 a32311a <=( a32310a  and  a32305a );
 a32315a <=( A234  and  A232 );
 a32316a <=( A203  and  a32315a );
 a32320a <=( A269  and  A266 );
 a32321a <=( (not A265)  and  a32320a );
 a32322a <=( a32321a  and  a32316a );
 a32326a <=( A167  and  (not A168) );
 a32327a <=( (not A169)  and  a32326a );
 a32331a <=( (not A200)  and  A199 );
 a32332a <=( A166  and  a32331a );
 a32333a <=( a32332a  and  a32327a );
 a32337a <=( A234  and  A232 );
 a32338a <=( A203  and  a32337a );
 a32342a <=( A269  and  (not A266) );
 a32343a <=( A265  and  a32342a );
 a32344a <=( a32343a  and  a32338a );
 a32348a <=( A167  and  (not A168) );
 a32349a <=( (not A169)  and  a32348a );
 a32353a <=( (not A200)  and  A199 );
 a32354a <=( A166  and  a32353a );
 a32355a <=( a32354a  and  a32349a );
 a32359a <=( A234  and  A233 );
 a32360a <=( A203  and  a32359a );
 a32364a <=( A302  and  (not A299) );
 a32365a <=( A298  and  a32364a );
 a32366a <=( a32365a  and  a32360a );
 a32370a <=( A167  and  (not A168) );
 a32371a <=( (not A169)  and  a32370a );
 a32375a <=( (not A200)  and  A199 );
 a32376a <=( A166  and  a32375a );
 a32377a <=( a32376a  and  a32371a );
 a32381a <=( A234  and  A233 );
 a32382a <=( A203  and  a32381a );
 a32386a <=( A302  and  A299 );
 a32387a <=( (not A298)  and  a32386a );
 a32388a <=( a32387a  and  a32382a );
 a32392a <=( A167  and  (not A168) );
 a32393a <=( (not A169)  and  a32392a );
 a32397a <=( (not A200)  and  A199 );
 a32398a <=( A166  and  a32397a );
 a32399a <=( a32398a  and  a32393a );
 a32403a <=( A234  and  A233 );
 a32404a <=( A203  and  a32403a );
 a32408a <=( A269  and  A266 );
 a32409a <=( (not A265)  and  a32408a );
 a32410a <=( a32409a  and  a32404a );
 a32414a <=( A167  and  (not A168) );
 a32415a <=( (not A169)  and  a32414a );
 a32419a <=( (not A200)  and  A199 );
 a32420a <=( A166  and  a32419a );
 a32421a <=( a32420a  and  a32415a );
 a32425a <=( A234  and  A233 );
 a32426a <=( A203  and  a32425a );
 a32430a <=( A269  and  (not A266) );
 a32431a <=( A265  and  a32430a );
 a32432a <=( a32431a  and  a32426a );
 a32436a <=( A167  and  (not A168) );
 a32437a <=( (not A169)  and  a32436a );
 a32441a <=( (not A200)  and  A199 );
 a32442a <=( A166  and  a32441a );
 a32443a <=( a32442a  and  a32437a );
 a32447a <=( A233  and  (not A232) );
 a32448a <=( A203  and  a32447a );
 a32452a <=( A300  and  A299 );
 a32453a <=( A236  and  a32452a );
 a32454a <=( a32453a  and  a32448a );
 a32458a <=( A167  and  (not A168) );
 a32459a <=( (not A169)  and  a32458a );
 a32463a <=( (not A200)  and  A199 );
 a32464a <=( A166  and  a32463a );
 a32465a <=( a32464a  and  a32459a );
 a32469a <=( A233  and  (not A232) );
 a32470a <=( A203  and  a32469a );
 a32474a <=( A300  and  A298 );
 a32475a <=( A236  and  a32474a );
 a32476a <=( a32475a  and  a32470a );
 a32480a <=( A167  and  (not A168) );
 a32481a <=( (not A169)  and  a32480a );
 a32485a <=( (not A200)  and  A199 );
 a32486a <=( A166  and  a32485a );
 a32487a <=( a32486a  and  a32481a );
 a32491a <=( A233  and  (not A232) );
 a32492a <=( A203  and  a32491a );
 a32496a <=( A267  and  A265 );
 a32497a <=( A236  and  a32496a );
 a32498a <=( a32497a  and  a32492a );
 a32502a <=( A167  and  (not A168) );
 a32503a <=( (not A169)  and  a32502a );
 a32507a <=( (not A200)  and  A199 );
 a32508a <=( A166  and  a32507a );
 a32509a <=( a32508a  and  a32503a );
 a32513a <=( A233  and  (not A232) );
 a32514a <=( A203  and  a32513a );
 a32518a <=( A267  and  A266 );
 a32519a <=( A236  and  a32518a );
 a32520a <=( a32519a  and  a32514a );
 a32524a <=( A167  and  (not A168) );
 a32525a <=( (not A169)  and  a32524a );
 a32529a <=( (not A200)  and  A199 );
 a32530a <=( A166  and  a32529a );
 a32531a <=( a32530a  and  a32525a );
 a32535a <=( (not A233)  and  A232 );
 a32536a <=( A203  and  a32535a );
 a32540a <=( A300  and  A299 );
 a32541a <=( A236  and  a32540a );
 a32542a <=( a32541a  and  a32536a );
 a32546a <=( A167  and  (not A168) );
 a32547a <=( (not A169)  and  a32546a );
 a32551a <=( (not A200)  and  A199 );
 a32552a <=( A166  and  a32551a );
 a32553a <=( a32552a  and  a32547a );
 a32557a <=( (not A233)  and  A232 );
 a32558a <=( A203  and  a32557a );
 a32562a <=( A300  and  A298 );
 a32563a <=( A236  and  a32562a );
 a32564a <=( a32563a  and  a32558a );
 a32568a <=( A167  and  (not A168) );
 a32569a <=( (not A169)  and  a32568a );
 a32573a <=( (not A200)  and  A199 );
 a32574a <=( A166  and  a32573a );
 a32575a <=( a32574a  and  a32569a );
 a32579a <=( (not A233)  and  A232 );
 a32580a <=( A203  and  a32579a );
 a32584a <=( A267  and  A265 );
 a32585a <=( A236  and  a32584a );
 a32586a <=( a32585a  and  a32580a );
 a32590a <=( A167  and  (not A168) );
 a32591a <=( (not A169)  and  a32590a );
 a32595a <=( (not A200)  and  A199 );
 a32596a <=( A166  and  a32595a );
 a32597a <=( a32596a  and  a32591a );
 a32601a <=( (not A233)  and  A232 );
 a32602a <=( A203  and  a32601a );
 a32606a <=( A267  and  A266 );
 a32607a <=( A236  and  a32606a );
 a32608a <=( a32607a  and  a32602a );
 a32612a <=( (not A168)  and  (not A169) );
 a32613a <=( (not A170)  and  a32612a );
 a32617a <=( A203  and  A200 );
 a32618a <=( (not A199)  and  a32617a );
 a32619a <=( a32618a  and  a32613a );
 a32623a <=( A236  and  A233 );
 a32624a <=( (not A232)  and  a32623a );
 a32628a <=( A302  and  (not A299) );
 a32629a <=( A298  and  a32628a );
 a32630a <=( a32629a  and  a32624a );
 a32634a <=( (not A168)  and  (not A169) );
 a32635a <=( (not A170)  and  a32634a );
 a32639a <=( A203  and  A200 );
 a32640a <=( (not A199)  and  a32639a );
 a32641a <=( a32640a  and  a32635a );
 a32645a <=( A236  and  A233 );
 a32646a <=( (not A232)  and  a32645a );
 a32650a <=( A302  and  A299 );
 a32651a <=( (not A298)  and  a32650a );
 a32652a <=( a32651a  and  a32646a );
 a32656a <=( (not A168)  and  (not A169) );
 a32657a <=( (not A170)  and  a32656a );
 a32661a <=( A203  and  A200 );
 a32662a <=( (not A199)  and  a32661a );
 a32663a <=( a32662a  and  a32657a );
 a32667a <=( A236  and  A233 );
 a32668a <=( (not A232)  and  a32667a );
 a32672a <=( A269  and  A266 );
 a32673a <=( (not A265)  and  a32672a );
 a32674a <=( a32673a  and  a32668a );
 a32678a <=( (not A168)  and  (not A169) );
 a32679a <=( (not A170)  and  a32678a );
 a32683a <=( A203  and  A200 );
 a32684a <=( (not A199)  and  a32683a );
 a32685a <=( a32684a  and  a32679a );
 a32689a <=( A236  and  A233 );
 a32690a <=( (not A232)  and  a32689a );
 a32694a <=( A269  and  (not A266) );
 a32695a <=( A265  and  a32694a );
 a32696a <=( a32695a  and  a32690a );
 a32700a <=( (not A168)  and  (not A169) );
 a32701a <=( (not A170)  and  a32700a );
 a32705a <=( A203  and  A200 );
 a32706a <=( (not A199)  and  a32705a );
 a32707a <=( a32706a  and  a32701a );
 a32711a <=( A236  and  (not A233) );
 a32712a <=( A232  and  a32711a );
 a32716a <=( A302  and  (not A299) );
 a32717a <=( A298  and  a32716a );
 a32718a <=( a32717a  and  a32712a );
 a32722a <=( (not A168)  and  (not A169) );
 a32723a <=( (not A170)  and  a32722a );
 a32727a <=( A203  and  A200 );
 a32728a <=( (not A199)  and  a32727a );
 a32729a <=( a32728a  and  a32723a );
 a32733a <=( A236  and  (not A233) );
 a32734a <=( A232  and  a32733a );
 a32738a <=( A302  and  A299 );
 a32739a <=( (not A298)  and  a32738a );
 a32740a <=( a32739a  and  a32734a );
 a32744a <=( (not A168)  and  (not A169) );
 a32745a <=( (not A170)  and  a32744a );
 a32749a <=( A203  and  A200 );
 a32750a <=( (not A199)  and  a32749a );
 a32751a <=( a32750a  and  a32745a );
 a32755a <=( A236  and  (not A233) );
 a32756a <=( A232  and  a32755a );
 a32760a <=( A269  and  A266 );
 a32761a <=( (not A265)  and  a32760a );
 a32762a <=( a32761a  and  a32756a );
 a32766a <=( (not A168)  and  (not A169) );
 a32767a <=( (not A170)  and  a32766a );
 a32771a <=( A203  and  A200 );
 a32772a <=( (not A199)  and  a32771a );
 a32773a <=( a32772a  and  a32767a );
 a32777a <=( A236  and  (not A233) );
 a32778a <=( A232  and  a32777a );
 a32782a <=( A269  and  (not A266) );
 a32783a <=( A265  and  a32782a );
 a32784a <=( a32783a  and  a32778a );
 a32788a <=( (not A168)  and  (not A169) );
 a32789a <=( (not A170)  and  a32788a );
 a32793a <=( A203  and  (not A200) );
 a32794a <=( A199  and  a32793a );
 a32795a <=( a32794a  and  a32789a );
 a32799a <=( A236  and  A233 );
 a32800a <=( (not A232)  and  a32799a );
 a32804a <=( A302  and  (not A299) );
 a32805a <=( A298  and  a32804a );
 a32806a <=( a32805a  and  a32800a );
 a32810a <=( (not A168)  and  (not A169) );
 a32811a <=( (not A170)  and  a32810a );
 a32815a <=( A203  and  (not A200) );
 a32816a <=( A199  and  a32815a );
 a32817a <=( a32816a  and  a32811a );
 a32821a <=( A236  and  A233 );
 a32822a <=( (not A232)  and  a32821a );
 a32826a <=( A302  and  A299 );
 a32827a <=( (not A298)  and  a32826a );
 a32828a <=( a32827a  and  a32822a );
 a32832a <=( (not A168)  and  (not A169) );
 a32833a <=( (not A170)  and  a32832a );
 a32837a <=( A203  and  (not A200) );
 a32838a <=( A199  and  a32837a );
 a32839a <=( a32838a  and  a32833a );
 a32843a <=( A236  and  A233 );
 a32844a <=( (not A232)  and  a32843a );
 a32848a <=( A269  and  A266 );
 a32849a <=( (not A265)  and  a32848a );
 a32850a <=( a32849a  and  a32844a );
 a32854a <=( (not A168)  and  (not A169) );
 a32855a <=( (not A170)  and  a32854a );
 a32859a <=( A203  and  (not A200) );
 a32860a <=( A199  and  a32859a );
 a32861a <=( a32860a  and  a32855a );
 a32865a <=( A236  and  A233 );
 a32866a <=( (not A232)  and  a32865a );
 a32870a <=( A269  and  (not A266) );
 a32871a <=( A265  and  a32870a );
 a32872a <=( a32871a  and  a32866a );
 a32876a <=( (not A168)  and  (not A169) );
 a32877a <=( (not A170)  and  a32876a );
 a32881a <=( A203  and  (not A200) );
 a32882a <=( A199  and  a32881a );
 a32883a <=( a32882a  and  a32877a );
 a32887a <=( A236  and  (not A233) );
 a32888a <=( A232  and  a32887a );
 a32892a <=( A302  and  (not A299) );
 a32893a <=( A298  and  a32892a );
 a32894a <=( a32893a  and  a32888a );
 a32898a <=( (not A168)  and  (not A169) );
 a32899a <=( (not A170)  and  a32898a );
 a32903a <=( A203  and  (not A200) );
 a32904a <=( A199  and  a32903a );
 a32905a <=( a32904a  and  a32899a );
 a32909a <=( A236  and  (not A233) );
 a32910a <=( A232  and  a32909a );
 a32914a <=( A302  and  A299 );
 a32915a <=( (not A298)  and  a32914a );
 a32916a <=( a32915a  and  a32910a );
 a32920a <=( (not A168)  and  (not A169) );
 a32921a <=( (not A170)  and  a32920a );
 a32925a <=( A203  and  (not A200) );
 a32926a <=( A199  and  a32925a );
 a32927a <=( a32926a  and  a32921a );
 a32931a <=( A236  and  (not A233) );
 a32932a <=( A232  and  a32931a );
 a32936a <=( A269  and  A266 );
 a32937a <=( (not A265)  and  a32936a );
 a32938a <=( a32937a  and  a32932a );
 a32942a <=( (not A168)  and  (not A169) );
 a32943a <=( (not A170)  and  a32942a );
 a32947a <=( A203  and  (not A200) );
 a32948a <=( A199  and  a32947a );
 a32949a <=( a32948a  and  a32943a );
 a32953a <=( A236  and  (not A233) );
 a32954a <=( A232  and  a32953a );
 a32958a <=( A269  and  (not A266) );
 a32959a <=( A265  and  a32958a );
 a32960a <=( a32959a  and  a32954a );
 a32964a <=( (not A166)  and  A167 );
 a32965a <=( A170  and  a32964a );
 a32969a <=( (not A201)  and  A200 );
 a32970a <=( A199  and  a32969a );
 a32971a <=( a32970a  and  a32965a );
 a32975a <=( A233  and  (not A232) );
 a32976a <=( (not A202)  and  a32975a );
 a32979a <=( A298  and  A236 );
 a32982a <=( A302  and  (not A299) );
 a32983a <=( a32982a  and  a32979a );
 a32984a <=( a32983a  and  a32976a );
 a32988a <=( (not A166)  and  A167 );
 a32989a <=( A170  and  a32988a );
 a32993a <=( (not A201)  and  A200 );
 a32994a <=( A199  and  a32993a );
 a32995a <=( a32994a  and  a32989a );
 a32999a <=( A233  and  (not A232) );
 a33000a <=( (not A202)  and  a32999a );
 a33003a <=( (not A298)  and  A236 );
 a33006a <=( A302  and  A299 );
 a33007a <=( a33006a  and  a33003a );
 a33008a <=( a33007a  and  a33000a );
 a33012a <=( (not A166)  and  A167 );
 a33013a <=( A170  and  a33012a );
 a33017a <=( (not A201)  and  A200 );
 a33018a <=( A199  and  a33017a );
 a33019a <=( a33018a  and  a33013a );
 a33023a <=( A233  and  (not A232) );
 a33024a <=( (not A202)  and  a33023a );
 a33027a <=( (not A265)  and  A236 );
 a33030a <=( A269  and  A266 );
 a33031a <=( a33030a  and  a33027a );
 a33032a <=( a33031a  and  a33024a );
 a33036a <=( (not A166)  and  A167 );
 a33037a <=( A170  and  a33036a );
 a33041a <=( (not A201)  and  A200 );
 a33042a <=( A199  and  a33041a );
 a33043a <=( a33042a  and  a33037a );
 a33047a <=( A233  and  (not A232) );
 a33048a <=( (not A202)  and  a33047a );
 a33051a <=( A265  and  A236 );
 a33054a <=( A269  and  (not A266) );
 a33055a <=( a33054a  and  a33051a );
 a33056a <=( a33055a  and  a33048a );
 a33060a <=( (not A166)  and  A167 );
 a33061a <=( A170  and  a33060a );
 a33065a <=( (not A201)  and  A200 );
 a33066a <=( A199  and  a33065a );
 a33067a <=( a33066a  and  a33061a );
 a33071a <=( (not A233)  and  A232 );
 a33072a <=( (not A202)  and  a33071a );
 a33075a <=( A298  and  A236 );
 a33078a <=( A302  and  (not A299) );
 a33079a <=( a33078a  and  a33075a );
 a33080a <=( a33079a  and  a33072a );
 a33084a <=( (not A166)  and  A167 );
 a33085a <=( A170  and  a33084a );
 a33089a <=( (not A201)  and  A200 );
 a33090a <=( A199  and  a33089a );
 a33091a <=( a33090a  and  a33085a );
 a33095a <=( (not A233)  and  A232 );
 a33096a <=( (not A202)  and  a33095a );
 a33099a <=( (not A298)  and  A236 );
 a33102a <=( A302  and  A299 );
 a33103a <=( a33102a  and  a33099a );
 a33104a <=( a33103a  and  a33096a );
 a33108a <=( (not A166)  and  A167 );
 a33109a <=( A170  and  a33108a );
 a33113a <=( (not A201)  and  A200 );
 a33114a <=( A199  and  a33113a );
 a33115a <=( a33114a  and  a33109a );
 a33119a <=( (not A233)  and  A232 );
 a33120a <=( (not A202)  and  a33119a );
 a33123a <=( (not A265)  and  A236 );
 a33126a <=( A269  and  A266 );
 a33127a <=( a33126a  and  a33123a );
 a33128a <=( a33127a  and  a33120a );
 a33132a <=( (not A166)  and  A167 );
 a33133a <=( A170  and  a33132a );
 a33137a <=( (not A201)  and  A200 );
 a33138a <=( A199  and  a33137a );
 a33139a <=( a33138a  and  a33133a );
 a33143a <=( (not A233)  and  A232 );
 a33144a <=( (not A202)  and  a33143a );
 a33147a <=( A265  and  A236 );
 a33150a <=( A269  and  (not A266) );
 a33151a <=( a33150a  and  a33147a );
 a33152a <=( a33151a  and  a33144a );
 a33156a <=( A166  and  (not A167) );
 a33157a <=( A170  and  a33156a );
 a33161a <=( (not A201)  and  A200 );
 a33162a <=( A199  and  a33161a );
 a33163a <=( a33162a  and  a33157a );
 a33167a <=( A233  and  (not A232) );
 a33168a <=( (not A202)  and  a33167a );
 a33171a <=( A298  and  A236 );
 a33174a <=( A302  and  (not A299) );
 a33175a <=( a33174a  and  a33171a );
 a33176a <=( a33175a  and  a33168a );
 a33180a <=( A166  and  (not A167) );
 a33181a <=( A170  and  a33180a );
 a33185a <=( (not A201)  and  A200 );
 a33186a <=( A199  and  a33185a );
 a33187a <=( a33186a  and  a33181a );
 a33191a <=( A233  and  (not A232) );
 a33192a <=( (not A202)  and  a33191a );
 a33195a <=( (not A298)  and  A236 );
 a33198a <=( A302  and  A299 );
 a33199a <=( a33198a  and  a33195a );
 a33200a <=( a33199a  and  a33192a );
 a33204a <=( A166  and  (not A167) );
 a33205a <=( A170  and  a33204a );
 a33209a <=( (not A201)  and  A200 );
 a33210a <=( A199  and  a33209a );
 a33211a <=( a33210a  and  a33205a );
 a33215a <=( A233  and  (not A232) );
 a33216a <=( (not A202)  and  a33215a );
 a33219a <=( (not A265)  and  A236 );
 a33222a <=( A269  and  A266 );
 a33223a <=( a33222a  and  a33219a );
 a33224a <=( a33223a  and  a33216a );
 a33228a <=( A166  and  (not A167) );
 a33229a <=( A170  and  a33228a );
 a33233a <=( (not A201)  and  A200 );
 a33234a <=( A199  and  a33233a );
 a33235a <=( a33234a  and  a33229a );
 a33239a <=( A233  and  (not A232) );
 a33240a <=( (not A202)  and  a33239a );
 a33243a <=( A265  and  A236 );
 a33246a <=( A269  and  (not A266) );
 a33247a <=( a33246a  and  a33243a );
 a33248a <=( a33247a  and  a33240a );
 a33252a <=( A166  and  (not A167) );
 a33253a <=( A170  and  a33252a );
 a33257a <=( (not A201)  and  A200 );
 a33258a <=( A199  and  a33257a );
 a33259a <=( a33258a  and  a33253a );
 a33263a <=( (not A233)  and  A232 );
 a33264a <=( (not A202)  and  a33263a );
 a33267a <=( A298  and  A236 );
 a33270a <=( A302  and  (not A299) );
 a33271a <=( a33270a  and  a33267a );
 a33272a <=( a33271a  and  a33264a );
 a33276a <=( A166  and  (not A167) );
 a33277a <=( A170  and  a33276a );
 a33281a <=( (not A201)  and  A200 );
 a33282a <=( A199  and  a33281a );
 a33283a <=( a33282a  and  a33277a );
 a33287a <=( (not A233)  and  A232 );
 a33288a <=( (not A202)  and  a33287a );
 a33291a <=( (not A298)  and  A236 );
 a33294a <=( A302  and  A299 );
 a33295a <=( a33294a  and  a33291a );
 a33296a <=( a33295a  and  a33288a );
 a33300a <=( A166  and  (not A167) );
 a33301a <=( A170  and  a33300a );
 a33305a <=( (not A201)  and  A200 );
 a33306a <=( A199  and  a33305a );
 a33307a <=( a33306a  and  a33301a );
 a33311a <=( (not A233)  and  A232 );
 a33312a <=( (not A202)  and  a33311a );
 a33315a <=( (not A265)  and  A236 );
 a33318a <=( A269  and  A266 );
 a33319a <=( a33318a  and  a33315a );
 a33320a <=( a33319a  and  a33312a );
 a33324a <=( A166  and  (not A167) );
 a33325a <=( A170  and  a33324a );
 a33329a <=( (not A201)  and  A200 );
 a33330a <=( A199  and  a33329a );
 a33331a <=( a33330a  and  a33325a );
 a33335a <=( (not A233)  and  A232 );
 a33336a <=( (not A202)  and  a33335a );
 a33339a <=( A265  and  A236 );
 a33342a <=( A269  and  (not A266) );
 a33343a <=( a33342a  and  a33339a );
 a33344a <=( a33343a  and  a33336a );
 a33348a <=( (not A202)  and  (not A201) );
 a33349a <=( A169  and  a33348a );
 a33353a <=( (not A235)  and  (not A234) );
 a33354a <=( (not A203)  and  a33353a );
 a33355a <=( a33354a  and  a33349a );
 a33359a <=( (not A268)  and  (not A267) );
 a33360a <=( (not A236)  and  a33359a );
 a33363a <=( (not A300)  and  (not A269) );
 a33366a <=( (not A302)  and  (not A301) );
 a33367a <=( a33366a  and  a33363a );
 a33368a <=( a33367a  and  a33360a );
 a33372a <=( (not A202)  and  (not A201) );
 a33373a <=( A169  and  a33372a );
 a33377a <=( (not A235)  and  (not A234) );
 a33378a <=( (not A203)  and  a33377a );
 a33379a <=( a33378a  and  a33373a );
 a33383a <=( (not A268)  and  (not A267) );
 a33384a <=( (not A236)  and  a33383a );
 a33387a <=( (not A298)  and  (not A269) );
 a33390a <=( (not A301)  and  (not A299) );
 a33391a <=( a33390a  and  a33387a );
 a33392a <=( a33391a  and  a33384a );
 a33396a <=( (not A202)  and  (not A201) );
 a33397a <=( A169  and  a33396a );
 a33401a <=( (not A235)  and  (not A234) );
 a33402a <=( (not A203)  and  a33401a );
 a33403a <=( a33402a  and  a33397a );
 a33407a <=( (not A266)  and  (not A265) );
 a33408a <=( (not A236)  and  a33407a );
 a33411a <=( (not A300)  and  (not A268) );
 a33414a <=( (not A302)  and  (not A301) );
 a33415a <=( a33414a  and  a33411a );
 a33416a <=( a33415a  and  a33408a );
 a33420a <=( (not A202)  and  (not A201) );
 a33421a <=( A169  and  a33420a );
 a33425a <=( (not A235)  and  (not A234) );
 a33426a <=( (not A203)  and  a33425a );
 a33427a <=( a33426a  and  a33421a );
 a33431a <=( (not A266)  and  (not A265) );
 a33432a <=( (not A236)  and  a33431a );
 a33435a <=( (not A298)  and  (not A268) );
 a33438a <=( (not A301)  and  (not A299) );
 a33439a <=( a33438a  and  a33435a );
 a33440a <=( a33439a  and  a33432a );
 a33444a <=( (not A202)  and  (not A201) );
 a33445a <=( A169  and  a33444a );
 a33449a <=( (not A233)  and  (not A232) );
 a33450a <=( (not A203)  and  a33449a );
 a33451a <=( a33450a  and  a33445a );
 a33455a <=( (not A268)  and  (not A267) );
 a33456a <=( (not A235)  and  a33455a );
 a33459a <=( (not A300)  and  (not A269) );
 a33462a <=( (not A302)  and  (not A301) );
 a33463a <=( a33462a  and  a33459a );
 a33464a <=( a33463a  and  a33456a );
 a33468a <=( (not A202)  and  (not A201) );
 a33469a <=( A169  and  a33468a );
 a33473a <=( (not A233)  and  (not A232) );
 a33474a <=( (not A203)  and  a33473a );
 a33475a <=( a33474a  and  a33469a );
 a33479a <=( (not A268)  and  (not A267) );
 a33480a <=( (not A235)  and  a33479a );
 a33483a <=( (not A298)  and  (not A269) );
 a33486a <=( (not A301)  and  (not A299) );
 a33487a <=( a33486a  and  a33483a );
 a33488a <=( a33487a  and  a33480a );
 a33492a <=( (not A202)  and  (not A201) );
 a33493a <=( A169  and  a33492a );
 a33497a <=( (not A233)  and  (not A232) );
 a33498a <=( (not A203)  and  a33497a );
 a33499a <=( a33498a  and  a33493a );
 a33503a <=( (not A266)  and  (not A265) );
 a33504a <=( (not A235)  and  a33503a );
 a33507a <=( (not A300)  and  (not A268) );
 a33510a <=( (not A302)  and  (not A301) );
 a33511a <=( a33510a  and  a33507a );
 a33512a <=( a33511a  and  a33504a );
 a33516a <=( (not A202)  and  (not A201) );
 a33517a <=( A169  and  a33516a );
 a33521a <=( (not A233)  and  (not A232) );
 a33522a <=( (not A203)  and  a33521a );
 a33523a <=( a33522a  and  a33517a );
 a33527a <=( (not A266)  and  (not A265) );
 a33528a <=( (not A235)  and  a33527a );
 a33531a <=( (not A298)  and  (not A268) );
 a33534a <=( (not A301)  and  (not A299) );
 a33535a <=( a33534a  and  a33531a );
 a33536a <=( a33535a  and  a33528a );
 a33540a <=( (not A200)  and  (not A199) );
 a33541a <=( A169  and  a33540a );
 a33545a <=( (not A235)  and  (not A234) );
 a33546a <=( (not A202)  and  a33545a );
 a33547a <=( a33546a  and  a33541a );
 a33551a <=( (not A268)  and  (not A267) );
 a33552a <=( (not A236)  and  a33551a );
 a33555a <=( (not A300)  and  (not A269) );
 a33558a <=( (not A302)  and  (not A301) );
 a33559a <=( a33558a  and  a33555a );
 a33560a <=( a33559a  and  a33552a );
 a33564a <=( (not A200)  and  (not A199) );
 a33565a <=( A169  and  a33564a );
 a33569a <=( (not A235)  and  (not A234) );
 a33570a <=( (not A202)  and  a33569a );
 a33571a <=( a33570a  and  a33565a );
 a33575a <=( (not A268)  and  (not A267) );
 a33576a <=( (not A236)  and  a33575a );
 a33579a <=( (not A298)  and  (not A269) );
 a33582a <=( (not A301)  and  (not A299) );
 a33583a <=( a33582a  and  a33579a );
 a33584a <=( a33583a  and  a33576a );
 a33588a <=( (not A200)  and  (not A199) );
 a33589a <=( A169  and  a33588a );
 a33593a <=( (not A235)  and  (not A234) );
 a33594a <=( (not A202)  and  a33593a );
 a33595a <=( a33594a  and  a33589a );
 a33599a <=( (not A266)  and  (not A265) );
 a33600a <=( (not A236)  and  a33599a );
 a33603a <=( (not A300)  and  (not A268) );
 a33606a <=( (not A302)  and  (not A301) );
 a33607a <=( a33606a  and  a33603a );
 a33608a <=( a33607a  and  a33600a );
 a33612a <=( (not A200)  and  (not A199) );
 a33613a <=( A169  and  a33612a );
 a33617a <=( (not A235)  and  (not A234) );
 a33618a <=( (not A202)  and  a33617a );
 a33619a <=( a33618a  and  a33613a );
 a33623a <=( (not A266)  and  (not A265) );
 a33624a <=( (not A236)  and  a33623a );
 a33627a <=( (not A298)  and  (not A268) );
 a33630a <=( (not A301)  and  (not A299) );
 a33631a <=( a33630a  and  a33627a );
 a33632a <=( a33631a  and  a33624a );
 a33636a <=( (not A200)  and  (not A199) );
 a33637a <=( A169  and  a33636a );
 a33641a <=( (not A233)  and  (not A232) );
 a33642a <=( (not A202)  and  a33641a );
 a33643a <=( a33642a  and  a33637a );
 a33647a <=( (not A268)  and  (not A267) );
 a33648a <=( (not A235)  and  a33647a );
 a33651a <=( (not A300)  and  (not A269) );
 a33654a <=( (not A302)  and  (not A301) );
 a33655a <=( a33654a  and  a33651a );
 a33656a <=( a33655a  and  a33648a );
 a33660a <=( (not A200)  and  (not A199) );
 a33661a <=( A169  and  a33660a );
 a33665a <=( (not A233)  and  (not A232) );
 a33666a <=( (not A202)  and  a33665a );
 a33667a <=( a33666a  and  a33661a );
 a33671a <=( (not A268)  and  (not A267) );
 a33672a <=( (not A235)  and  a33671a );
 a33675a <=( (not A298)  and  (not A269) );
 a33678a <=( (not A301)  and  (not A299) );
 a33679a <=( a33678a  and  a33675a );
 a33680a <=( a33679a  and  a33672a );
 a33684a <=( (not A200)  and  (not A199) );
 a33685a <=( A169  and  a33684a );
 a33689a <=( (not A233)  and  (not A232) );
 a33690a <=( (not A202)  and  a33689a );
 a33691a <=( a33690a  and  a33685a );
 a33695a <=( (not A266)  and  (not A265) );
 a33696a <=( (not A235)  and  a33695a );
 a33699a <=( (not A300)  and  (not A268) );
 a33702a <=( (not A302)  and  (not A301) );
 a33703a <=( a33702a  and  a33699a );
 a33704a <=( a33703a  and  a33696a );
 a33708a <=( (not A200)  and  (not A199) );
 a33709a <=( A169  and  a33708a );
 a33713a <=( (not A233)  and  (not A232) );
 a33714a <=( (not A202)  and  a33713a );
 a33715a <=( a33714a  and  a33709a );
 a33719a <=( (not A266)  and  (not A265) );
 a33720a <=( (not A235)  and  a33719a );
 a33723a <=( (not A298)  and  (not A268) );
 a33726a <=( (not A301)  and  (not A299) );
 a33727a <=( a33726a  and  a33723a );
 a33728a <=( a33727a  and  a33720a );
 a33732a <=( (not A166)  and  (not A167) );
 a33733a <=( (not A169)  and  a33732a );
 a33737a <=( (not A235)  and  (not A234) );
 a33738a <=( A202  and  a33737a );
 a33739a <=( a33738a  and  a33733a );
 a33743a <=( (not A268)  and  (not A267) );
 a33744a <=( (not A236)  and  a33743a );
 a33747a <=( (not A300)  and  (not A269) );
 a33750a <=( (not A302)  and  (not A301) );
 a33751a <=( a33750a  and  a33747a );
 a33752a <=( a33751a  and  a33744a );
 a33756a <=( (not A166)  and  (not A167) );
 a33757a <=( (not A169)  and  a33756a );
 a33761a <=( (not A235)  and  (not A234) );
 a33762a <=( A202  and  a33761a );
 a33763a <=( a33762a  and  a33757a );
 a33767a <=( (not A268)  and  (not A267) );
 a33768a <=( (not A236)  and  a33767a );
 a33771a <=( (not A298)  and  (not A269) );
 a33774a <=( (not A301)  and  (not A299) );
 a33775a <=( a33774a  and  a33771a );
 a33776a <=( a33775a  and  a33768a );
 a33780a <=( (not A166)  and  (not A167) );
 a33781a <=( (not A169)  and  a33780a );
 a33785a <=( (not A235)  and  (not A234) );
 a33786a <=( A202  and  a33785a );
 a33787a <=( a33786a  and  a33781a );
 a33791a <=( (not A266)  and  (not A265) );
 a33792a <=( (not A236)  and  a33791a );
 a33795a <=( (not A300)  and  (not A268) );
 a33798a <=( (not A302)  and  (not A301) );
 a33799a <=( a33798a  and  a33795a );
 a33800a <=( a33799a  and  a33792a );
 a33804a <=( (not A166)  and  (not A167) );
 a33805a <=( (not A169)  and  a33804a );
 a33809a <=( (not A235)  and  (not A234) );
 a33810a <=( A202  and  a33809a );
 a33811a <=( a33810a  and  a33805a );
 a33815a <=( (not A266)  and  (not A265) );
 a33816a <=( (not A236)  and  a33815a );
 a33819a <=( (not A298)  and  (not A268) );
 a33822a <=( (not A301)  and  (not A299) );
 a33823a <=( a33822a  and  a33819a );
 a33824a <=( a33823a  and  a33816a );
 a33828a <=( (not A166)  and  (not A167) );
 a33829a <=( (not A169)  and  a33828a );
 a33833a <=( (not A233)  and  (not A232) );
 a33834a <=( A202  and  a33833a );
 a33835a <=( a33834a  and  a33829a );
 a33839a <=( (not A268)  and  (not A267) );
 a33840a <=( (not A235)  and  a33839a );
 a33843a <=( (not A300)  and  (not A269) );
 a33846a <=( (not A302)  and  (not A301) );
 a33847a <=( a33846a  and  a33843a );
 a33848a <=( a33847a  and  a33840a );
 a33852a <=( (not A166)  and  (not A167) );
 a33853a <=( (not A169)  and  a33852a );
 a33857a <=( (not A233)  and  (not A232) );
 a33858a <=( A202  and  a33857a );
 a33859a <=( a33858a  and  a33853a );
 a33863a <=( (not A268)  and  (not A267) );
 a33864a <=( (not A235)  and  a33863a );
 a33867a <=( (not A298)  and  (not A269) );
 a33870a <=( (not A301)  and  (not A299) );
 a33871a <=( a33870a  and  a33867a );
 a33872a <=( a33871a  and  a33864a );
 a33876a <=( (not A166)  and  (not A167) );
 a33877a <=( (not A169)  and  a33876a );
 a33881a <=( (not A233)  and  (not A232) );
 a33882a <=( A202  and  a33881a );
 a33883a <=( a33882a  and  a33877a );
 a33887a <=( (not A266)  and  (not A265) );
 a33888a <=( (not A235)  and  a33887a );
 a33891a <=( (not A300)  and  (not A268) );
 a33894a <=( (not A302)  and  (not A301) );
 a33895a <=( a33894a  and  a33891a );
 a33896a <=( a33895a  and  a33888a );
 a33900a <=( (not A166)  and  (not A167) );
 a33901a <=( (not A169)  and  a33900a );
 a33905a <=( (not A233)  and  (not A232) );
 a33906a <=( A202  and  a33905a );
 a33907a <=( a33906a  and  a33901a );
 a33911a <=( (not A266)  and  (not A265) );
 a33912a <=( (not A235)  and  a33911a );
 a33915a <=( (not A298)  and  (not A268) );
 a33918a <=( (not A301)  and  (not A299) );
 a33919a <=( a33918a  and  a33915a );
 a33920a <=( a33919a  and  a33912a );
 a33924a <=( A167  and  (not A168) );
 a33925a <=( (not A169)  and  a33924a );
 a33929a <=( A200  and  (not A199) );
 a33930a <=( A166  and  a33929a );
 a33931a <=( a33930a  and  a33925a );
 a33935a <=( A233  and  (not A232) );
 a33936a <=( A203  and  a33935a );
 a33939a <=( A298  and  A236 );
 a33942a <=( A302  and  (not A299) );
 a33943a <=( a33942a  and  a33939a );
 a33944a <=( a33943a  and  a33936a );
 a33948a <=( A167  and  (not A168) );
 a33949a <=( (not A169)  and  a33948a );
 a33953a <=( A200  and  (not A199) );
 a33954a <=( A166  and  a33953a );
 a33955a <=( a33954a  and  a33949a );
 a33959a <=( A233  and  (not A232) );
 a33960a <=( A203  and  a33959a );
 a33963a <=( (not A298)  and  A236 );
 a33966a <=( A302  and  A299 );
 a33967a <=( a33966a  and  a33963a );
 a33968a <=( a33967a  and  a33960a );
 a33972a <=( A167  and  (not A168) );
 a33973a <=( (not A169)  and  a33972a );
 a33977a <=( A200  and  (not A199) );
 a33978a <=( A166  and  a33977a );
 a33979a <=( a33978a  and  a33973a );
 a33983a <=( A233  and  (not A232) );
 a33984a <=( A203  and  a33983a );
 a33987a <=( (not A265)  and  A236 );
 a33990a <=( A269  and  A266 );
 a33991a <=( a33990a  and  a33987a );
 a33992a <=( a33991a  and  a33984a );
 a33996a <=( A167  and  (not A168) );
 a33997a <=( (not A169)  and  a33996a );
 a34001a <=( A200  and  (not A199) );
 a34002a <=( A166  and  a34001a );
 a34003a <=( a34002a  and  a33997a );
 a34007a <=( A233  and  (not A232) );
 a34008a <=( A203  and  a34007a );
 a34011a <=( A265  and  A236 );
 a34014a <=( A269  and  (not A266) );
 a34015a <=( a34014a  and  a34011a );
 a34016a <=( a34015a  and  a34008a );
 a34020a <=( A167  and  (not A168) );
 a34021a <=( (not A169)  and  a34020a );
 a34025a <=( A200  and  (not A199) );
 a34026a <=( A166  and  a34025a );
 a34027a <=( a34026a  and  a34021a );
 a34031a <=( (not A233)  and  A232 );
 a34032a <=( A203  and  a34031a );
 a34035a <=( A298  and  A236 );
 a34038a <=( A302  and  (not A299) );
 a34039a <=( a34038a  and  a34035a );
 a34040a <=( a34039a  and  a34032a );
 a34044a <=( A167  and  (not A168) );
 a34045a <=( (not A169)  and  a34044a );
 a34049a <=( A200  and  (not A199) );
 a34050a <=( A166  and  a34049a );
 a34051a <=( a34050a  and  a34045a );
 a34055a <=( (not A233)  and  A232 );
 a34056a <=( A203  and  a34055a );
 a34059a <=( (not A298)  and  A236 );
 a34062a <=( A302  and  A299 );
 a34063a <=( a34062a  and  a34059a );
 a34064a <=( a34063a  and  a34056a );
 a34068a <=( A167  and  (not A168) );
 a34069a <=( (not A169)  and  a34068a );
 a34073a <=( A200  and  (not A199) );
 a34074a <=( A166  and  a34073a );
 a34075a <=( a34074a  and  a34069a );
 a34079a <=( (not A233)  and  A232 );
 a34080a <=( A203  and  a34079a );
 a34083a <=( (not A265)  and  A236 );
 a34086a <=( A269  and  A266 );
 a34087a <=( a34086a  and  a34083a );
 a34088a <=( a34087a  and  a34080a );
 a34092a <=( A167  and  (not A168) );
 a34093a <=( (not A169)  and  a34092a );
 a34097a <=( A200  and  (not A199) );
 a34098a <=( A166  and  a34097a );
 a34099a <=( a34098a  and  a34093a );
 a34103a <=( (not A233)  and  A232 );
 a34104a <=( A203  and  a34103a );
 a34107a <=( A265  and  A236 );
 a34110a <=( A269  and  (not A266) );
 a34111a <=( a34110a  and  a34107a );
 a34112a <=( a34111a  and  a34104a );
 a34116a <=( A167  and  (not A168) );
 a34117a <=( (not A169)  and  a34116a );
 a34121a <=( (not A200)  and  A199 );
 a34122a <=( A166  and  a34121a );
 a34123a <=( a34122a  and  a34117a );
 a34127a <=( A233  and  (not A232) );
 a34128a <=( A203  and  a34127a );
 a34131a <=( A298  and  A236 );
 a34134a <=( A302  and  (not A299) );
 a34135a <=( a34134a  and  a34131a );
 a34136a <=( a34135a  and  a34128a );
 a34140a <=( A167  and  (not A168) );
 a34141a <=( (not A169)  and  a34140a );
 a34145a <=( (not A200)  and  A199 );
 a34146a <=( A166  and  a34145a );
 a34147a <=( a34146a  and  a34141a );
 a34151a <=( A233  and  (not A232) );
 a34152a <=( A203  and  a34151a );
 a34155a <=( (not A298)  and  A236 );
 a34158a <=( A302  and  A299 );
 a34159a <=( a34158a  and  a34155a );
 a34160a <=( a34159a  and  a34152a );
 a34164a <=( A167  and  (not A168) );
 a34165a <=( (not A169)  and  a34164a );
 a34169a <=( (not A200)  and  A199 );
 a34170a <=( A166  and  a34169a );
 a34171a <=( a34170a  and  a34165a );
 a34175a <=( A233  and  (not A232) );
 a34176a <=( A203  and  a34175a );
 a34179a <=( (not A265)  and  A236 );
 a34182a <=( A269  and  A266 );
 a34183a <=( a34182a  and  a34179a );
 a34184a <=( a34183a  and  a34176a );
 a34188a <=( A167  and  (not A168) );
 a34189a <=( (not A169)  and  a34188a );
 a34193a <=( (not A200)  and  A199 );
 a34194a <=( A166  and  a34193a );
 a34195a <=( a34194a  and  a34189a );
 a34199a <=( A233  and  (not A232) );
 a34200a <=( A203  and  a34199a );
 a34203a <=( A265  and  A236 );
 a34206a <=( A269  and  (not A266) );
 a34207a <=( a34206a  and  a34203a );
 a34208a <=( a34207a  and  a34200a );
 a34212a <=( A167  and  (not A168) );
 a34213a <=( (not A169)  and  a34212a );
 a34217a <=( (not A200)  and  A199 );
 a34218a <=( A166  and  a34217a );
 a34219a <=( a34218a  and  a34213a );
 a34223a <=( (not A233)  and  A232 );
 a34224a <=( A203  and  a34223a );
 a34227a <=( A298  and  A236 );
 a34230a <=( A302  and  (not A299) );
 a34231a <=( a34230a  and  a34227a );
 a34232a <=( a34231a  and  a34224a );
 a34236a <=( A167  and  (not A168) );
 a34237a <=( (not A169)  and  a34236a );
 a34241a <=( (not A200)  and  A199 );
 a34242a <=( A166  and  a34241a );
 a34243a <=( a34242a  and  a34237a );
 a34247a <=( (not A233)  and  A232 );
 a34248a <=( A203  and  a34247a );
 a34251a <=( (not A298)  and  A236 );
 a34254a <=( A302  and  A299 );
 a34255a <=( a34254a  and  a34251a );
 a34256a <=( a34255a  and  a34248a );
 a34260a <=( A167  and  (not A168) );
 a34261a <=( (not A169)  and  a34260a );
 a34265a <=( (not A200)  and  A199 );
 a34266a <=( A166  and  a34265a );
 a34267a <=( a34266a  and  a34261a );
 a34271a <=( (not A233)  and  A232 );
 a34272a <=( A203  and  a34271a );
 a34275a <=( (not A265)  and  A236 );
 a34278a <=( A269  and  A266 );
 a34279a <=( a34278a  and  a34275a );
 a34280a <=( a34279a  and  a34272a );
 a34284a <=( A167  and  (not A168) );
 a34285a <=( (not A169)  and  a34284a );
 a34289a <=( (not A200)  and  A199 );
 a34290a <=( A166  and  a34289a );
 a34291a <=( a34290a  and  a34285a );
 a34295a <=( (not A233)  and  A232 );
 a34296a <=( A203  and  a34295a );
 a34299a <=( A265  and  A236 );
 a34302a <=( A269  and  (not A266) );
 a34303a <=( a34302a  and  a34299a );
 a34304a <=( a34303a  and  a34296a );
 a34308a <=( (not A168)  and  (not A169) );
 a34309a <=( (not A170)  and  a34308a );
 a34313a <=( (not A235)  and  (not A234) );
 a34314a <=( A202  and  a34313a );
 a34315a <=( a34314a  and  a34309a );
 a34319a <=( (not A268)  and  (not A267) );
 a34320a <=( (not A236)  and  a34319a );
 a34323a <=( (not A300)  and  (not A269) );
 a34326a <=( (not A302)  and  (not A301) );
 a34327a <=( a34326a  and  a34323a );
 a34328a <=( a34327a  and  a34320a );
 a34332a <=( (not A168)  and  (not A169) );
 a34333a <=( (not A170)  and  a34332a );
 a34337a <=( (not A235)  and  (not A234) );
 a34338a <=( A202  and  a34337a );
 a34339a <=( a34338a  and  a34333a );
 a34343a <=( (not A268)  and  (not A267) );
 a34344a <=( (not A236)  and  a34343a );
 a34347a <=( (not A298)  and  (not A269) );
 a34350a <=( (not A301)  and  (not A299) );
 a34351a <=( a34350a  and  a34347a );
 a34352a <=( a34351a  and  a34344a );
 a34356a <=( (not A168)  and  (not A169) );
 a34357a <=( (not A170)  and  a34356a );
 a34361a <=( (not A235)  and  (not A234) );
 a34362a <=( A202  and  a34361a );
 a34363a <=( a34362a  and  a34357a );
 a34367a <=( (not A266)  and  (not A265) );
 a34368a <=( (not A236)  and  a34367a );
 a34371a <=( (not A300)  and  (not A268) );
 a34374a <=( (not A302)  and  (not A301) );
 a34375a <=( a34374a  and  a34371a );
 a34376a <=( a34375a  and  a34368a );
 a34380a <=( (not A168)  and  (not A169) );
 a34381a <=( (not A170)  and  a34380a );
 a34385a <=( (not A235)  and  (not A234) );
 a34386a <=( A202  and  a34385a );
 a34387a <=( a34386a  and  a34381a );
 a34391a <=( (not A266)  and  (not A265) );
 a34392a <=( (not A236)  and  a34391a );
 a34395a <=( (not A298)  and  (not A268) );
 a34398a <=( (not A301)  and  (not A299) );
 a34399a <=( a34398a  and  a34395a );
 a34400a <=( a34399a  and  a34392a );
 a34404a <=( (not A168)  and  (not A169) );
 a34405a <=( (not A170)  and  a34404a );
 a34409a <=( (not A233)  and  (not A232) );
 a34410a <=( A202  and  a34409a );
 a34411a <=( a34410a  and  a34405a );
 a34415a <=( (not A268)  and  (not A267) );
 a34416a <=( (not A235)  and  a34415a );
 a34419a <=( (not A300)  and  (not A269) );
 a34422a <=( (not A302)  and  (not A301) );
 a34423a <=( a34422a  and  a34419a );
 a34424a <=( a34423a  and  a34416a );
 a34428a <=( (not A168)  and  (not A169) );
 a34429a <=( (not A170)  and  a34428a );
 a34433a <=( (not A233)  and  (not A232) );
 a34434a <=( A202  and  a34433a );
 a34435a <=( a34434a  and  a34429a );
 a34439a <=( (not A268)  and  (not A267) );
 a34440a <=( (not A235)  and  a34439a );
 a34443a <=( (not A298)  and  (not A269) );
 a34446a <=( (not A301)  and  (not A299) );
 a34447a <=( a34446a  and  a34443a );
 a34448a <=( a34447a  and  a34440a );
 a34452a <=( (not A168)  and  (not A169) );
 a34453a <=( (not A170)  and  a34452a );
 a34457a <=( (not A233)  and  (not A232) );
 a34458a <=( A202  and  a34457a );
 a34459a <=( a34458a  and  a34453a );
 a34463a <=( (not A266)  and  (not A265) );
 a34464a <=( (not A235)  and  a34463a );
 a34467a <=( (not A300)  and  (not A268) );
 a34470a <=( (not A302)  and  (not A301) );
 a34471a <=( a34470a  and  a34467a );
 a34472a <=( a34471a  and  a34464a );
 a34476a <=( (not A168)  and  (not A169) );
 a34477a <=( (not A170)  and  a34476a );
 a34481a <=( (not A233)  and  (not A232) );
 a34482a <=( A202  and  a34481a );
 a34483a <=( a34482a  and  a34477a );
 a34487a <=( (not A266)  and  (not A265) );
 a34488a <=( (not A235)  and  a34487a );
 a34491a <=( (not A298)  and  (not A268) );
 a34494a <=( (not A301)  and  (not A299) );
 a34495a <=( a34494a  and  a34491a );
 a34496a <=( a34495a  and  a34488a );
 a34500a <=( (not A201)  and  A166 );
 a34501a <=( A168  and  a34500a );
 a34504a <=( (not A203)  and  (not A202) );
 a34507a <=( (not A235)  and  (not A234) );
 a34508a <=( a34507a  and  a34504a );
 a34509a <=( a34508a  and  a34501a );
 a34513a <=( (not A268)  and  (not A267) );
 a34514a <=( (not A236)  and  a34513a );
 a34517a <=( (not A300)  and  (not A269) );
 a34520a <=( (not A302)  and  (not A301) );
 a34521a <=( a34520a  and  a34517a );
 a34522a <=( a34521a  and  a34514a );
 a34526a <=( (not A201)  and  A166 );
 a34527a <=( A168  and  a34526a );
 a34530a <=( (not A203)  and  (not A202) );
 a34533a <=( (not A235)  and  (not A234) );
 a34534a <=( a34533a  and  a34530a );
 a34535a <=( a34534a  and  a34527a );
 a34539a <=( (not A268)  and  (not A267) );
 a34540a <=( (not A236)  and  a34539a );
 a34543a <=( (not A298)  and  (not A269) );
 a34546a <=( (not A301)  and  (not A299) );
 a34547a <=( a34546a  and  a34543a );
 a34548a <=( a34547a  and  a34540a );
 a34552a <=( (not A201)  and  A166 );
 a34553a <=( A168  and  a34552a );
 a34556a <=( (not A203)  and  (not A202) );
 a34559a <=( (not A235)  and  (not A234) );
 a34560a <=( a34559a  and  a34556a );
 a34561a <=( a34560a  and  a34553a );
 a34565a <=( (not A266)  and  (not A265) );
 a34566a <=( (not A236)  and  a34565a );
 a34569a <=( (not A300)  and  (not A268) );
 a34572a <=( (not A302)  and  (not A301) );
 a34573a <=( a34572a  and  a34569a );
 a34574a <=( a34573a  and  a34566a );
 a34578a <=( (not A201)  and  A166 );
 a34579a <=( A168  and  a34578a );
 a34582a <=( (not A203)  and  (not A202) );
 a34585a <=( (not A235)  and  (not A234) );
 a34586a <=( a34585a  and  a34582a );
 a34587a <=( a34586a  and  a34579a );
 a34591a <=( (not A266)  and  (not A265) );
 a34592a <=( (not A236)  and  a34591a );
 a34595a <=( (not A298)  and  (not A268) );
 a34598a <=( (not A301)  and  (not A299) );
 a34599a <=( a34598a  and  a34595a );
 a34600a <=( a34599a  and  a34592a );
 a34604a <=( (not A201)  and  A166 );
 a34605a <=( A168  and  a34604a );
 a34608a <=( (not A203)  and  (not A202) );
 a34611a <=( (not A233)  and  (not A232) );
 a34612a <=( a34611a  and  a34608a );
 a34613a <=( a34612a  and  a34605a );
 a34617a <=( (not A268)  and  (not A267) );
 a34618a <=( (not A235)  and  a34617a );
 a34621a <=( (not A300)  and  (not A269) );
 a34624a <=( (not A302)  and  (not A301) );
 a34625a <=( a34624a  and  a34621a );
 a34626a <=( a34625a  and  a34618a );
 a34630a <=( (not A201)  and  A166 );
 a34631a <=( A168  and  a34630a );
 a34634a <=( (not A203)  and  (not A202) );
 a34637a <=( (not A233)  and  (not A232) );
 a34638a <=( a34637a  and  a34634a );
 a34639a <=( a34638a  and  a34631a );
 a34643a <=( (not A268)  and  (not A267) );
 a34644a <=( (not A235)  and  a34643a );
 a34647a <=( (not A298)  and  (not A269) );
 a34650a <=( (not A301)  and  (not A299) );
 a34651a <=( a34650a  and  a34647a );
 a34652a <=( a34651a  and  a34644a );
 a34656a <=( (not A201)  and  A166 );
 a34657a <=( A168  and  a34656a );
 a34660a <=( (not A203)  and  (not A202) );
 a34663a <=( (not A233)  and  (not A232) );
 a34664a <=( a34663a  and  a34660a );
 a34665a <=( a34664a  and  a34657a );
 a34669a <=( (not A266)  and  (not A265) );
 a34670a <=( (not A235)  and  a34669a );
 a34673a <=( (not A300)  and  (not A268) );
 a34676a <=( (not A302)  and  (not A301) );
 a34677a <=( a34676a  and  a34673a );
 a34678a <=( a34677a  and  a34670a );
 a34682a <=( (not A201)  and  A166 );
 a34683a <=( A168  and  a34682a );
 a34686a <=( (not A203)  and  (not A202) );
 a34689a <=( (not A233)  and  (not A232) );
 a34690a <=( a34689a  and  a34686a );
 a34691a <=( a34690a  and  a34683a );
 a34695a <=( (not A266)  and  (not A265) );
 a34696a <=( (not A235)  and  a34695a );
 a34699a <=( (not A298)  and  (not A268) );
 a34702a <=( (not A301)  and  (not A299) );
 a34703a <=( a34702a  and  a34699a );
 a34704a <=( a34703a  and  a34696a );
 a34708a <=( (not A199)  and  A166 );
 a34709a <=( A168  and  a34708a );
 a34712a <=( (not A202)  and  (not A200) );
 a34715a <=( (not A235)  and  (not A234) );
 a34716a <=( a34715a  and  a34712a );
 a34717a <=( a34716a  and  a34709a );
 a34721a <=( (not A268)  and  (not A267) );
 a34722a <=( (not A236)  and  a34721a );
 a34725a <=( (not A300)  and  (not A269) );
 a34728a <=( (not A302)  and  (not A301) );
 a34729a <=( a34728a  and  a34725a );
 a34730a <=( a34729a  and  a34722a );
 a34734a <=( (not A199)  and  A166 );
 a34735a <=( A168  and  a34734a );
 a34738a <=( (not A202)  and  (not A200) );
 a34741a <=( (not A235)  and  (not A234) );
 a34742a <=( a34741a  and  a34738a );
 a34743a <=( a34742a  and  a34735a );
 a34747a <=( (not A268)  and  (not A267) );
 a34748a <=( (not A236)  and  a34747a );
 a34751a <=( (not A298)  and  (not A269) );
 a34754a <=( (not A301)  and  (not A299) );
 a34755a <=( a34754a  and  a34751a );
 a34756a <=( a34755a  and  a34748a );
 a34760a <=( (not A199)  and  A166 );
 a34761a <=( A168  and  a34760a );
 a34764a <=( (not A202)  and  (not A200) );
 a34767a <=( (not A235)  and  (not A234) );
 a34768a <=( a34767a  and  a34764a );
 a34769a <=( a34768a  and  a34761a );
 a34773a <=( (not A266)  and  (not A265) );
 a34774a <=( (not A236)  and  a34773a );
 a34777a <=( (not A300)  and  (not A268) );
 a34780a <=( (not A302)  and  (not A301) );
 a34781a <=( a34780a  and  a34777a );
 a34782a <=( a34781a  and  a34774a );
 a34786a <=( (not A199)  and  A166 );
 a34787a <=( A168  and  a34786a );
 a34790a <=( (not A202)  and  (not A200) );
 a34793a <=( (not A235)  and  (not A234) );
 a34794a <=( a34793a  and  a34790a );
 a34795a <=( a34794a  and  a34787a );
 a34799a <=( (not A266)  and  (not A265) );
 a34800a <=( (not A236)  and  a34799a );
 a34803a <=( (not A298)  and  (not A268) );
 a34806a <=( (not A301)  and  (not A299) );
 a34807a <=( a34806a  and  a34803a );
 a34808a <=( a34807a  and  a34800a );
 a34812a <=( (not A199)  and  A166 );
 a34813a <=( A168  and  a34812a );
 a34816a <=( (not A202)  and  (not A200) );
 a34819a <=( (not A233)  and  (not A232) );
 a34820a <=( a34819a  and  a34816a );
 a34821a <=( a34820a  and  a34813a );
 a34825a <=( (not A268)  and  (not A267) );
 a34826a <=( (not A235)  and  a34825a );
 a34829a <=( (not A300)  and  (not A269) );
 a34832a <=( (not A302)  and  (not A301) );
 a34833a <=( a34832a  and  a34829a );
 a34834a <=( a34833a  and  a34826a );
 a34838a <=( (not A199)  and  A166 );
 a34839a <=( A168  and  a34838a );
 a34842a <=( (not A202)  and  (not A200) );
 a34845a <=( (not A233)  and  (not A232) );
 a34846a <=( a34845a  and  a34842a );
 a34847a <=( a34846a  and  a34839a );
 a34851a <=( (not A268)  and  (not A267) );
 a34852a <=( (not A235)  and  a34851a );
 a34855a <=( (not A298)  and  (not A269) );
 a34858a <=( (not A301)  and  (not A299) );
 a34859a <=( a34858a  and  a34855a );
 a34860a <=( a34859a  and  a34852a );
 a34864a <=( (not A199)  and  A166 );
 a34865a <=( A168  and  a34864a );
 a34868a <=( (not A202)  and  (not A200) );
 a34871a <=( (not A233)  and  (not A232) );
 a34872a <=( a34871a  and  a34868a );
 a34873a <=( a34872a  and  a34865a );
 a34877a <=( (not A266)  and  (not A265) );
 a34878a <=( (not A235)  and  a34877a );
 a34881a <=( (not A300)  and  (not A268) );
 a34884a <=( (not A302)  and  (not A301) );
 a34885a <=( a34884a  and  a34881a );
 a34886a <=( a34885a  and  a34878a );
 a34890a <=( (not A199)  and  A166 );
 a34891a <=( A168  and  a34890a );
 a34894a <=( (not A202)  and  (not A200) );
 a34897a <=( (not A233)  and  (not A232) );
 a34898a <=( a34897a  and  a34894a );
 a34899a <=( a34898a  and  a34891a );
 a34903a <=( (not A266)  and  (not A265) );
 a34904a <=( (not A235)  and  a34903a );
 a34907a <=( (not A298)  and  (not A268) );
 a34910a <=( (not A301)  and  (not A299) );
 a34911a <=( a34910a  and  a34907a );
 a34912a <=( a34911a  and  a34904a );
 a34916a <=( (not A201)  and  A167 );
 a34917a <=( A168  and  a34916a );
 a34920a <=( (not A203)  and  (not A202) );
 a34923a <=( (not A235)  and  (not A234) );
 a34924a <=( a34923a  and  a34920a );
 a34925a <=( a34924a  and  a34917a );
 a34929a <=( (not A268)  and  (not A267) );
 a34930a <=( (not A236)  and  a34929a );
 a34933a <=( (not A300)  and  (not A269) );
 a34936a <=( (not A302)  and  (not A301) );
 a34937a <=( a34936a  and  a34933a );
 a34938a <=( a34937a  and  a34930a );
 a34942a <=( (not A201)  and  A167 );
 a34943a <=( A168  and  a34942a );
 a34946a <=( (not A203)  and  (not A202) );
 a34949a <=( (not A235)  and  (not A234) );
 a34950a <=( a34949a  and  a34946a );
 a34951a <=( a34950a  and  a34943a );
 a34955a <=( (not A268)  and  (not A267) );
 a34956a <=( (not A236)  and  a34955a );
 a34959a <=( (not A298)  and  (not A269) );
 a34962a <=( (not A301)  and  (not A299) );
 a34963a <=( a34962a  and  a34959a );
 a34964a <=( a34963a  and  a34956a );
 a34968a <=( (not A201)  and  A167 );
 a34969a <=( A168  and  a34968a );
 a34972a <=( (not A203)  and  (not A202) );
 a34975a <=( (not A235)  and  (not A234) );
 a34976a <=( a34975a  and  a34972a );
 a34977a <=( a34976a  and  a34969a );
 a34981a <=( (not A266)  and  (not A265) );
 a34982a <=( (not A236)  and  a34981a );
 a34985a <=( (not A300)  and  (not A268) );
 a34988a <=( (not A302)  and  (not A301) );
 a34989a <=( a34988a  and  a34985a );
 a34990a <=( a34989a  and  a34982a );
 a34994a <=( (not A201)  and  A167 );
 a34995a <=( A168  and  a34994a );
 a34998a <=( (not A203)  and  (not A202) );
 a35001a <=( (not A235)  and  (not A234) );
 a35002a <=( a35001a  and  a34998a );
 a35003a <=( a35002a  and  a34995a );
 a35007a <=( (not A266)  and  (not A265) );
 a35008a <=( (not A236)  and  a35007a );
 a35011a <=( (not A298)  and  (not A268) );
 a35014a <=( (not A301)  and  (not A299) );
 a35015a <=( a35014a  and  a35011a );
 a35016a <=( a35015a  and  a35008a );
 a35020a <=( (not A201)  and  A167 );
 a35021a <=( A168  and  a35020a );
 a35024a <=( (not A203)  and  (not A202) );
 a35027a <=( (not A233)  and  (not A232) );
 a35028a <=( a35027a  and  a35024a );
 a35029a <=( a35028a  and  a35021a );
 a35033a <=( (not A268)  and  (not A267) );
 a35034a <=( (not A235)  and  a35033a );
 a35037a <=( (not A300)  and  (not A269) );
 a35040a <=( (not A302)  and  (not A301) );
 a35041a <=( a35040a  and  a35037a );
 a35042a <=( a35041a  and  a35034a );
 a35046a <=( (not A201)  and  A167 );
 a35047a <=( A168  and  a35046a );
 a35050a <=( (not A203)  and  (not A202) );
 a35053a <=( (not A233)  and  (not A232) );
 a35054a <=( a35053a  and  a35050a );
 a35055a <=( a35054a  and  a35047a );
 a35059a <=( (not A268)  and  (not A267) );
 a35060a <=( (not A235)  and  a35059a );
 a35063a <=( (not A298)  and  (not A269) );
 a35066a <=( (not A301)  and  (not A299) );
 a35067a <=( a35066a  and  a35063a );
 a35068a <=( a35067a  and  a35060a );
 a35072a <=( (not A201)  and  A167 );
 a35073a <=( A168  and  a35072a );
 a35076a <=( (not A203)  and  (not A202) );
 a35079a <=( (not A233)  and  (not A232) );
 a35080a <=( a35079a  and  a35076a );
 a35081a <=( a35080a  and  a35073a );
 a35085a <=( (not A266)  and  (not A265) );
 a35086a <=( (not A235)  and  a35085a );
 a35089a <=( (not A300)  and  (not A268) );
 a35092a <=( (not A302)  and  (not A301) );
 a35093a <=( a35092a  and  a35089a );
 a35094a <=( a35093a  and  a35086a );
 a35098a <=( (not A201)  and  A167 );
 a35099a <=( A168  and  a35098a );
 a35102a <=( (not A203)  and  (not A202) );
 a35105a <=( (not A233)  and  (not A232) );
 a35106a <=( a35105a  and  a35102a );
 a35107a <=( a35106a  and  a35099a );
 a35111a <=( (not A266)  and  (not A265) );
 a35112a <=( (not A235)  and  a35111a );
 a35115a <=( (not A298)  and  (not A268) );
 a35118a <=( (not A301)  and  (not A299) );
 a35119a <=( a35118a  and  a35115a );
 a35120a <=( a35119a  and  a35112a );
 a35124a <=( (not A199)  and  A167 );
 a35125a <=( A168  and  a35124a );
 a35128a <=( (not A202)  and  (not A200) );
 a35131a <=( (not A235)  and  (not A234) );
 a35132a <=( a35131a  and  a35128a );
 a35133a <=( a35132a  and  a35125a );
 a35137a <=( (not A268)  and  (not A267) );
 a35138a <=( (not A236)  and  a35137a );
 a35141a <=( (not A300)  and  (not A269) );
 a35144a <=( (not A302)  and  (not A301) );
 a35145a <=( a35144a  and  a35141a );
 a35146a <=( a35145a  and  a35138a );
 a35150a <=( (not A199)  and  A167 );
 a35151a <=( A168  and  a35150a );
 a35154a <=( (not A202)  and  (not A200) );
 a35157a <=( (not A235)  and  (not A234) );
 a35158a <=( a35157a  and  a35154a );
 a35159a <=( a35158a  and  a35151a );
 a35163a <=( (not A268)  and  (not A267) );
 a35164a <=( (not A236)  and  a35163a );
 a35167a <=( (not A298)  and  (not A269) );
 a35170a <=( (not A301)  and  (not A299) );
 a35171a <=( a35170a  and  a35167a );
 a35172a <=( a35171a  and  a35164a );
 a35176a <=( (not A199)  and  A167 );
 a35177a <=( A168  and  a35176a );
 a35180a <=( (not A202)  and  (not A200) );
 a35183a <=( (not A235)  and  (not A234) );
 a35184a <=( a35183a  and  a35180a );
 a35185a <=( a35184a  and  a35177a );
 a35189a <=( (not A266)  and  (not A265) );
 a35190a <=( (not A236)  and  a35189a );
 a35193a <=( (not A300)  and  (not A268) );
 a35196a <=( (not A302)  and  (not A301) );
 a35197a <=( a35196a  and  a35193a );
 a35198a <=( a35197a  and  a35190a );
 a35202a <=( (not A199)  and  A167 );
 a35203a <=( A168  and  a35202a );
 a35206a <=( (not A202)  and  (not A200) );
 a35209a <=( (not A235)  and  (not A234) );
 a35210a <=( a35209a  and  a35206a );
 a35211a <=( a35210a  and  a35203a );
 a35215a <=( (not A266)  and  (not A265) );
 a35216a <=( (not A236)  and  a35215a );
 a35219a <=( (not A298)  and  (not A268) );
 a35222a <=( (not A301)  and  (not A299) );
 a35223a <=( a35222a  and  a35219a );
 a35224a <=( a35223a  and  a35216a );
 a35228a <=( (not A199)  and  A167 );
 a35229a <=( A168  and  a35228a );
 a35232a <=( (not A202)  and  (not A200) );
 a35235a <=( (not A233)  and  (not A232) );
 a35236a <=( a35235a  and  a35232a );
 a35237a <=( a35236a  and  a35229a );
 a35241a <=( (not A268)  and  (not A267) );
 a35242a <=( (not A235)  and  a35241a );
 a35245a <=( (not A300)  and  (not A269) );
 a35248a <=( (not A302)  and  (not A301) );
 a35249a <=( a35248a  and  a35245a );
 a35250a <=( a35249a  and  a35242a );
 a35254a <=( (not A199)  and  A167 );
 a35255a <=( A168  and  a35254a );
 a35258a <=( (not A202)  and  (not A200) );
 a35261a <=( (not A233)  and  (not A232) );
 a35262a <=( a35261a  and  a35258a );
 a35263a <=( a35262a  and  a35255a );
 a35267a <=( (not A268)  and  (not A267) );
 a35268a <=( (not A235)  and  a35267a );
 a35271a <=( (not A298)  and  (not A269) );
 a35274a <=( (not A301)  and  (not A299) );
 a35275a <=( a35274a  and  a35271a );
 a35276a <=( a35275a  and  a35268a );
 a35280a <=( (not A199)  and  A167 );
 a35281a <=( A168  and  a35280a );
 a35284a <=( (not A202)  and  (not A200) );
 a35287a <=( (not A233)  and  (not A232) );
 a35288a <=( a35287a  and  a35284a );
 a35289a <=( a35288a  and  a35281a );
 a35293a <=( (not A266)  and  (not A265) );
 a35294a <=( (not A235)  and  a35293a );
 a35297a <=( (not A300)  and  (not A268) );
 a35300a <=( (not A302)  and  (not A301) );
 a35301a <=( a35300a  and  a35297a );
 a35302a <=( a35301a  and  a35294a );
 a35306a <=( (not A199)  and  A167 );
 a35307a <=( A168  and  a35306a );
 a35310a <=( (not A202)  and  (not A200) );
 a35313a <=( (not A233)  and  (not A232) );
 a35314a <=( a35313a  and  a35310a );
 a35315a <=( a35314a  and  a35307a );
 a35319a <=( (not A266)  and  (not A265) );
 a35320a <=( (not A235)  and  a35319a );
 a35323a <=( (not A298)  and  (not A268) );
 a35326a <=( (not A301)  and  (not A299) );
 a35327a <=( a35326a  and  a35323a );
 a35328a <=( a35327a  and  a35320a );
 a35332a <=( (not A202)  and  (not A201) );
 a35333a <=( A169  and  a35332a );
 a35336a <=( (not A234)  and  (not A203) );
 a35339a <=( (not A236)  and  (not A235) );
 a35340a <=( a35339a  and  a35336a );
 a35341a <=( a35340a  and  a35333a );
 a35345a <=( (not A269)  and  (not A268) );
 a35346a <=( (not A267)  and  a35345a );
 a35349a <=( A299  and  A298 );
 a35352a <=( (not A301)  and  (not A300) );
 a35353a <=( a35352a  and  a35349a );
 a35354a <=( a35353a  and  a35346a );
 a35358a <=( (not A202)  and  (not A201) );
 a35359a <=( A169  and  a35358a );
 a35362a <=( (not A234)  and  (not A203) );
 a35365a <=( (not A236)  and  (not A235) );
 a35366a <=( a35365a  and  a35362a );
 a35367a <=( a35366a  and  a35359a );
 a35371a <=( (not A267)  and  A266 );
 a35372a <=( A265  and  a35371a );
 a35375a <=( (not A300)  and  (not A268) );
 a35378a <=( (not A302)  and  (not A301) );
 a35379a <=( a35378a  and  a35375a );
 a35380a <=( a35379a  and  a35372a );
 a35384a <=( (not A202)  and  (not A201) );
 a35385a <=( A169  and  a35384a );
 a35388a <=( (not A234)  and  (not A203) );
 a35391a <=( (not A236)  and  (not A235) );
 a35392a <=( a35391a  and  a35388a );
 a35393a <=( a35392a  and  a35385a );
 a35397a <=( (not A267)  and  A266 );
 a35398a <=( A265  and  a35397a );
 a35401a <=( (not A298)  and  (not A268) );
 a35404a <=( (not A301)  and  (not A299) );
 a35405a <=( a35404a  and  a35401a );
 a35406a <=( a35405a  and  a35398a );
 a35410a <=( (not A202)  and  (not A201) );
 a35411a <=( A169  and  a35410a );
 a35414a <=( (not A234)  and  (not A203) );
 a35417a <=( (not A236)  and  (not A235) );
 a35418a <=( a35417a  and  a35414a );
 a35419a <=( a35418a  and  a35411a );
 a35423a <=( (not A268)  and  (not A266) );
 a35424a <=( (not A265)  and  a35423a );
 a35427a <=( A299  and  A298 );
 a35430a <=( (not A301)  and  (not A300) );
 a35431a <=( a35430a  and  a35427a );
 a35432a <=( a35431a  and  a35424a );
 a35436a <=( (not A202)  and  (not A201) );
 a35437a <=( A169  and  a35436a );
 a35440a <=( A232  and  (not A203) );
 a35443a <=( (not A234)  and  A233 );
 a35444a <=( a35443a  and  a35440a );
 a35445a <=( a35444a  and  a35437a );
 a35449a <=( (not A268)  and  (not A267) );
 a35450a <=( (not A235)  and  a35449a );
 a35453a <=( (not A300)  and  (not A269) );
 a35456a <=( (not A302)  and  (not A301) );
 a35457a <=( a35456a  and  a35453a );
 a35458a <=( a35457a  and  a35450a );
 a35462a <=( (not A202)  and  (not A201) );
 a35463a <=( A169  and  a35462a );
 a35466a <=( A232  and  (not A203) );
 a35469a <=( (not A234)  and  A233 );
 a35470a <=( a35469a  and  a35466a );
 a35471a <=( a35470a  and  a35463a );
 a35475a <=( (not A268)  and  (not A267) );
 a35476a <=( (not A235)  and  a35475a );
 a35479a <=( (not A298)  and  (not A269) );
 a35482a <=( (not A301)  and  (not A299) );
 a35483a <=( a35482a  and  a35479a );
 a35484a <=( a35483a  and  a35476a );
 a35488a <=( (not A202)  and  (not A201) );
 a35489a <=( A169  and  a35488a );
 a35492a <=( A232  and  (not A203) );
 a35495a <=( (not A234)  and  A233 );
 a35496a <=( a35495a  and  a35492a );
 a35497a <=( a35496a  and  a35489a );
 a35501a <=( (not A266)  and  (not A265) );
 a35502a <=( (not A235)  and  a35501a );
 a35505a <=( (not A300)  and  (not A268) );
 a35508a <=( (not A302)  and  (not A301) );
 a35509a <=( a35508a  and  a35505a );
 a35510a <=( a35509a  and  a35502a );
 a35514a <=( (not A202)  and  (not A201) );
 a35515a <=( A169  and  a35514a );
 a35518a <=( A232  and  (not A203) );
 a35521a <=( (not A234)  and  A233 );
 a35522a <=( a35521a  and  a35518a );
 a35523a <=( a35522a  and  a35515a );
 a35527a <=( (not A266)  and  (not A265) );
 a35528a <=( (not A235)  and  a35527a );
 a35531a <=( (not A298)  and  (not A268) );
 a35534a <=( (not A301)  and  (not A299) );
 a35535a <=( a35534a  and  a35531a );
 a35536a <=( a35535a  and  a35528a );
 a35540a <=( (not A202)  and  (not A201) );
 a35541a <=( A169  and  a35540a );
 a35544a <=( (not A232)  and  (not A203) );
 a35547a <=( (not A235)  and  (not A233) );
 a35548a <=( a35547a  and  a35544a );
 a35549a <=( a35548a  and  a35541a );
 a35553a <=( (not A269)  and  (not A268) );
 a35554a <=( (not A267)  and  a35553a );
 a35557a <=( A299  and  A298 );
 a35560a <=( (not A301)  and  (not A300) );
 a35561a <=( a35560a  and  a35557a );
 a35562a <=( a35561a  and  a35554a );
 a35566a <=( (not A202)  and  (not A201) );
 a35567a <=( A169  and  a35566a );
 a35570a <=( (not A232)  and  (not A203) );
 a35573a <=( (not A235)  and  (not A233) );
 a35574a <=( a35573a  and  a35570a );
 a35575a <=( a35574a  and  a35567a );
 a35579a <=( (not A267)  and  A266 );
 a35580a <=( A265  and  a35579a );
 a35583a <=( (not A300)  and  (not A268) );
 a35586a <=( (not A302)  and  (not A301) );
 a35587a <=( a35586a  and  a35583a );
 a35588a <=( a35587a  and  a35580a );
 a35592a <=( (not A202)  and  (not A201) );
 a35593a <=( A169  and  a35592a );
 a35596a <=( (not A232)  and  (not A203) );
 a35599a <=( (not A235)  and  (not A233) );
 a35600a <=( a35599a  and  a35596a );
 a35601a <=( a35600a  and  a35593a );
 a35605a <=( (not A267)  and  A266 );
 a35606a <=( A265  and  a35605a );
 a35609a <=( (not A298)  and  (not A268) );
 a35612a <=( (not A301)  and  (not A299) );
 a35613a <=( a35612a  and  a35609a );
 a35614a <=( a35613a  and  a35606a );
 a35618a <=( (not A202)  and  (not A201) );
 a35619a <=( A169  and  a35618a );
 a35622a <=( (not A232)  and  (not A203) );
 a35625a <=( (not A235)  and  (not A233) );
 a35626a <=( a35625a  and  a35622a );
 a35627a <=( a35626a  and  a35619a );
 a35631a <=( (not A268)  and  (not A266) );
 a35632a <=( (not A265)  and  a35631a );
 a35635a <=( A299  and  A298 );
 a35638a <=( (not A301)  and  (not A300) );
 a35639a <=( a35638a  and  a35635a );
 a35640a <=( a35639a  and  a35632a );
 a35644a <=( A200  and  A199 );
 a35645a <=( A169  and  a35644a );
 a35648a <=( (not A202)  and  (not A201) );
 a35651a <=( (not A235)  and  (not A234) );
 a35652a <=( a35651a  and  a35648a );
 a35653a <=( a35652a  and  a35645a );
 a35657a <=( (not A268)  and  (not A267) );
 a35658a <=( (not A236)  and  a35657a );
 a35661a <=( (not A300)  and  (not A269) );
 a35664a <=( (not A302)  and  (not A301) );
 a35665a <=( a35664a  and  a35661a );
 a35666a <=( a35665a  and  a35658a );
 a35670a <=( A200  and  A199 );
 a35671a <=( A169  and  a35670a );
 a35674a <=( (not A202)  and  (not A201) );
 a35677a <=( (not A235)  and  (not A234) );
 a35678a <=( a35677a  and  a35674a );
 a35679a <=( a35678a  and  a35671a );
 a35683a <=( (not A268)  and  (not A267) );
 a35684a <=( (not A236)  and  a35683a );
 a35687a <=( (not A298)  and  (not A269) );
 a35690a <=( (not A301)  and  (not A299) );
 a35691a <=( a35690a  and  a35687a );
 a35692a <=( a35691a  and  a35684a );
 a35696a <=( A200  and  A199 );
 a35697a <=( A169  and  a35696a );
 a35700a <=( (not A202)  and  (not A201) );
 a35703a <=( (not A235)  and  (not A234) );
 a35704a <=( a35703a  and  a35700a );
 a35705a <=( a35704a  and  a35697a );
 a35709a <=( (not A266)  and  (not A265) );
 a35710a <=( (not A236)  and  a35709a );
 a35713a <=( (not A300)  and  (not A268) );
 a35716a <=( (not A302)  and  (not A301) );
 a35717a <=( a35716a  and  a35713a );
 a35718a <=( a35717a  and  a35710a );
 a35722a <=( A200  and  A199 );
 a35723a <=( A169  and  a35722a );
 a35726a <=( (not A202)  and  (not A201) );
 a35729a <=( (not A235)  and  (not A234) );
 a35730a <=( a35729a  and  a35726a );
 a35731a <=( a35730a  and  a35723a );
 a35735a <=( (not A266)  and  (not A265) );
 a35736a <=( (not A236)  and  a35735a );
 a35739a <=( (not A298)  and  (not A268) );
 a35742a <=( (not A301)  and  (not A299) );
 a35743a <=( a35742a  and  a35739a );
 a35744a <=( a35743a  and  a35736a );
 a35748a <=( A200  and  A199 );
 a35749a <=( A169  and  a35748a );
 a35752a <=( (not A202)  and  (not A201) );
 a35755a <=( (not A233)  and  (not A232) );
 a35756a <=( a35755a  and  a35752a );
 a35757a <=( a35756a  and  a35749a );
 a35761a <=( (not A268)  and  (not A267) );
 a35762a <=( (not A235)  and  a35761a );
 a35765a <=( (not A300)  and  (not A269) );
 a35768a <=( (not A302)  and  (not A301) );
 a35769a <=( a35768a  and  a35765a );
 a35770a <=( a35769a  and  a35762a );
 a35774a <=( A200  and  A199 );
 a35775a <=( A169  and  a35774a );
 a35778a <=( (not A202)  and  (not A201) );
 a35781a <=( (not A233)  and  (not A232) );
 a35782a <=( a35781a  and  a35778a );
 a35783a <=( a35782a  and  a35775a );
 a35787a <=( (not A268)  and  (not A267) );
 a35788a <=( (not A235)  and  a35787a );
 a35791a <=( (not A298)  and  (not A269) );
 a35794a <=( (not A301)  and  (not A299) );
 a35795a <=( a35794a  and  a35791a );
 a35796a <=( a35795a  and  a35788a );
 a35800a <=( A200  and  A199 );
 a35801a <=( A169  and  a35800a );
 a35804a <=( (not A202)  and  (not A201) );
 a35807a <=( (not A233)  and  (not A232) );
 a35808a <=( a35807a  and  a35804a );
 a35809a <=( a35808a  and  a35801a );
 a35813a <=( (not A266)  and  (not A265) );
 a35814a <=( (not A235)  and  a35813a );
 a35817a <=( (not A300)  and  (not A268) );
 a35820a <=( (not A302)  and  (not A301) );
 a35821a <=( a35820a  and  a35817a );
 a35822a <=( a35821a  and  a35814a );
 a35826a <=( A200  and  A199 );
 a35827a <=( A169  and  a35826a );
 a35830a <=( (not A202)  and  (not A201) );
 a35833a <=( (not A233)  and  (not A232) );
 a35834a <=( a35833a  and  a35830a );
 a35835a <=( a35834a  and  a35827a );
 a35839a <=( (not A266)  and  (not A265) );
 a35840a <=( (not A235)  and  a35839a );
 a35843a <=( (not A298)  and  (not A268) );
 a35846a <=( (not A301)  and  (not A299) );
 a35847a <=( a35846a  and  a35843a );
 a35848a <=( a35847a  and  a35840a );
 a35852a <=( (not A200)  and  (not A199) );
 a35853a <=( A169  and  a35852a );
 a35856a <=( (not A234)  and  (not A202) );
 a35859a <=( (not A236)  and  (not A235) );
 a35860a <=( a35859a  and  a35856a );
 a35861a <=( a35860a  and  a35853a );
 a35865a <=( (not A269)  and  (not A268) );
 a35866a <=( (not A267)  and  a35865a );
 a35869a <=( A299  and  A298 );
 a35872a <=( (not A301)  and  (not A300) );
 a35873a <=( a35872a  and  a35869a );
 a35874a <=( a35873a  and  a35866a );
 a35878a <=( (not A200)  and  (not A199) );
 a35879a <=( A169  and  a35878a );
 a35882a <=( (not A234)  and  (not A202) );
 a35885a <=( (not A236)  and  (not A235) );
 a35886a <=( a35885a  and  a35882a );
 a35887a <=( a35886a  and  a35879a );
 a35891a <=( (not A267)  and  A266 );
 a35892a <=( A265  and  a35891a );
 a35895a <=( (not A300)  and  (not A268) );
 a35898a <=( (not A302)  and  (not A301) );
 a35899a <=( a35898a  and  a35895a );
 a35900a <=( a35899a  and  a35892a );
 a35904a <=( (not A200)  and  (not A199) );
 a35905a <=( A169  and  a35904a );
 a35908a <=( (not A234)  and  (not A202) );
 a35911a <=( (not A236)  and  (not A235) );
 a35912a <=( a35911a  and  a35908a );
 a35913a <=( a35912a  and  a35905a );
 a35917a <=( (not A267)  and  A266 );
 a35918a <=( A265  and  a35917a );
 a35921a <=( (not A298)  and  (not A268) );
 a35924a <=( (not A301)  and  (not A299) );
 a35925a <=( a35924a  and  a35921a );
 a35926a <=( a35925a  and  a35918a );
 a35930a <=( (not A200)  and  (not A199) );
 a35931a <=( A169  and  a35930a );
 a35934a <=( (not A234)  and  (not A202) );
 a35937a <=( (not A236)  and  (not A235) );
 a35938a <=( a35937a  and  a35934a );
 a35939a <=( a35938a  and  a35931a );
 a35943a <=( (not A268)  and  (not A266) );
 a35944a <=( (not A265)  and  a35943a );
 a35947a <=( A299  and  A298 );
 a35950a <=( (not A301)  and  (not A300) );
 a35951a <=( a35950a  and  a35947a );
 a35952a <=( a35951a  and  a35944a );
 a35956a <=( (not A200)  and  (not A199) );
 a35957a <=( A169  and  a35956a );
 a35960a <=( A232  and  (not A202) );
 a35963a <=( (not A234)  and  A233 );
 a35964a <=( a35963a  and  a35960a );
 a35965a <=( a35964a  and  a35957a );
 a35969a <=( (not A268)  and  (not A267) );
 a35970a <=( (not A235)  and  a35969a );
 a35973a <=( (not A300)  and  (not A269) );
 a35976a <=( (not A302)  and  (not A301) );
 a35977a <=( a35976a  and  a35973a );
 a35978a <=( a35977a  and  a35970a );
 a35982a <=( (not A200)  and  (not A199) );
 a35983a <=( A169  and  a35982a );
 a35986a <=( A232  and  (not A202) );
 a35989a <=( (not A234)  and  A233 );
 a35990a <=( a35989a  and  a35986a );
 a35991a <=( a35990a  and  a35983a );
 a35995a <=( (not A268)  and  (not A267) );
 a35996a <=( (not A235)  and  a35995a );
 a35999a <=( (not A298)  and  (not A269) );
 a36002a <=( (not A301)  and  (not A299) );
 a36003a <=( a36002a  and  a35999a );
 a36004a <=( a36003a  and  a35996a );
 a36008a <=( (not A200)  and  (not A199) );
 a36009a <=( A169  and  a36008a );
 a36012a <=( A232  and  (not A202) );
 a36015a <=( (not A234)  and  A233 );
 a36016a <=( a36015a  and  a36012a );
 a36017a <=( a36016a  and  a36009a );
 a36021a <=( (not A266)  and  (not A265) );
 a36022a <=( (not A235)  and  a36021a );
 a36025a <=( (not A300)  and  (not A268) );
 a36028a <=( (not A302)  and  (not A301) );
 a36029a <=( a36028a  and  a36025a );
 a36030a <=( a36029a  and  a36022a );
 a36034a <=( (not A200)  and  (not A199) );
 a36035a <=( A169  and  a36034a );
 a36038a <=( A232  and  (not A202) );
 a36041a <=( (not A234)  and  A233 );
 a36042a <=( a36041a  and  a36038a );
 a36043a <=( a36042a  and  a36035a );
 a36047a <=( (not A266)  and  (not A265) );
 a36048a <=( (not A235)  and  a36047a );
 a36051a <=( (not A298)  and  (not A268) );
 a36054a <=( (not A301)  and  (not A299) );
 a36055a <=( a36054a  and  a36051a );
 a36056a <=( a36055a  and  a36048a );
 a36060a <=( (not A200)  and  (not A199) );
 a36061a <=( A169  and  a36060a );
 a36064a <=( (not A232)  and  (not A202) );
 a36067a <=( (not A235)  and  (not A233) );
 a36068a <=( a36067a  and  a36064a );
 a36069a <=( a36068a  and  a36061a );
 a36073a <=( (not A269)  and  (not A268) );
 a36074a <=( (not A267)  and  a36073a );
 a36077a <=( A299  and  A298 );
 a36080a <=( (not A301)  and  (not A300) );
 a36081a <=( a36080a  and  a36077a );
 a36082a <=( a36081a  and  a36074a );
 a36086a <=( (not A200)  and  (not A199) );
 a36087a <=( A169  and  a36086a );
 a36090a <=( (not A232)  and  (not A202) );
 a36093a <=( (not A235)  and  (not A233) );
 a36094a <=( a36093a  and  a36090a );
 a36095a <=( a36094a  and  a36087a );
 a36099a <=( (not A267)  and  A266 );
 a36100a <=( A265  and  a36099a );
 a36103a <=( (not A300)  and  (not A268) );
 a36106a <=( (not A302)  and  (not A301) );
 a36107a <=( a36106a  and  a36103a );
 a36108a <=( a36107a  and  a36100a );
 a36112a <=( (not A200)  and  (not A199) );
 a36113a <=( A169  and  a36112a );
 a36116a <=( (not A232)  and  (not A202) );
 a36119a <=( (not A235)  and  (not A233) );
 a36120a <=( a36119a  and  a36116a );
 a36121a <=( a36120a  and  a36113a );
 a36125a <=( (not A267)  and  A266 );
 a36126a <=( A265  and  a36125a );
 a36129a <=( (not A298)  and  (not A268) );
 a36132a <=( (not A301)  and  (not A299) );
 a36133a <=( a36132a  and  a36129a );
 a36134a <=( a36133a  and  a36126a );
 a36138a <=( (not A200)  and  (not A199) );
 a36139a <=( A169  and  a36138a );
 a36142a <=( (not A232)  and  (not A202) );
 a36145a <=( (not A235)  and  (not A233) );
 a36146a <=( a36145a  and  a36142a );
 a36147a <=( a36146a  and  a36139a );
 a36151a <=( (not A268)  and  (not A266) );
 a36152a <=( (not A265)  and  a36151a );
 a36155a <=( A299  and  A298 );
 a36158a <=( (not A301)  and  (not A300) );
 a36159a <=( a36158a  and  a36155a );
 a36160a <=( a36159a  and  a36152a );
 a36164a <=( (not A166)  and  (not A167) );
 a36165a <=( (not A169)  and  a36164a );
 a36168a <=( (not A234)  and  A202 );
 a36171a <=( (not A236)  and  (not A235) );
 a36172a <=( a36171a  and  a36168a );
 a36173a <=( a36172a  and  a36165a );
 a36177a <=( (not A269)  and  (not A268) );
 a36178a <=( (not A267)  and  a36177a );
 a36181a <=( A299  and  A298 );
 a36184a <=( (not A301)  and  (not A300) );
 a36185a <=( a36184a  and  a36181a );
 a36186a <=( a36185a  and  a36178a );
 a36190a <=( (not A166)  and  (not A167) );
 a36191a <=( (not A169)  and  a36190a );
 a36194a <=( (not A234)  and  A202 );
 a36197a <=( (not A236)  and  (not A235) );
 a36198a <=( a36197a  and  a36194a );
 a36199a <=( a36198a  and  a36191a );
 a36203a <=( (not A267)  and  A266 );
 a36204a <=( A265  and  a36203a );
 a36207a <=( (not A300)  and  (not A268) );
 a36210a <=( (not A302)  and  (not A301) );
 a36211a <=( a36210a  and  a36207a );
 a36212a <=( a36211a  and  a36204a );
 a36216a <=( (not A166)  and  (not A167) );
 a36217a <=( (not A169)  and  a36216a );
 a36220a <=( (not A234)  and  A202 );
 a36223a <=( (not A236)  and  (not A235) );
 a36224a <=( a36223a  and  a36220a );
 a36225a <=( a36224a  and  a36217a );
 a36229a <=( (not A267)  and  A266 );
 a36230a <=( A265  and  a36229a );
 a36233a <=( (not A298)  and  (not A268) );
 a36236a <=( (not A301)  and  (not A299) );
 a36237a <=( a36236a  and  a36233a );
 a36238a <=( a36237a  and  a36230a );
 a36242a <=( (not A166)  and  (not A167) );
 a36243a <=( (not A169)  and  a36242a );
 a36246a <=( (not A234)  and  A202 );
 a36249a <=( (not A236)  and  (not A235) );
 a36250a <=( a36249a  and  a36246a );
 a36251a <=( a36250a  and  a36243a );
 a36255a <=( (not A268)  and  (not A266) );
 a36256a <=( (not A265)  and  a36255a );
 a36259a <=( A299  and  A298 );
 a36262a <=( (not A301)  and  (not A300) );
 a36263a <=( a36262a  and  a36259a );
 a36264a <=( a36263a  and  a36256a );
 a36268a <=( (not A166)  and  (not A167) );
 a36269a <=( (not A169)  and  a36268a );
 a36272a <=( A232  and  A202 );
 a36275a <=( (not A234)  and  A233 );
 a36276a <=( a36275a  and  a36272a );
 a36277a <=( a36276a  and  a36269a );
 a36281a <=( (not A268)  and  (not A267) );
 a36282a <=( (not A235)  and  a36281a );
 a36285a <=( (not A300)  and  (not A269) );
 a36288a <=( (not A302)  and  (not A301) );
 a36289a <=( a36288a  and  a36285a );
 a36290a <=( a36289a  and  a36282a );
 a36294a <=( (not A166)  and  (not A167) );
 a36295a <=( (not A169)  and  a36294a );
 a36298a <=( A232  and  A202 );
 a36301a <=( (not A234)  and  A233 );
 a36302a <=( a36301a  and  a36298a );
 a36303a <=( a36302a  and  a36295a );
 a36307a <=( (not A268)  and  (not A267) );
 a36308a <=( (not A235)  and  a36307a );
 a36311a <=( (not A298)  and  (not A269) );
 a36314a <=( (not A301)  and  (not A299) );
 a36315a <=( a36314a  and  a36311a );
 a36316a <=( a36315a  and  a36308a );
 a36320a <=( (not A166)  and  (not A167) );
 a36321a <=( (not A169)  and  a36320a );
 a36324a <=( A232  and  A202 );
 a36327a <=( (not A234)  and  A233 );
 a36328a <=( a36327a  and  a36324a );
 a36329a <=( a36328a  and  a36321a );
 a36333a <=( (not A266)  and  (not A265) );
 a36334a <=( (not A235)  and  a36333a );
 a36337a <=( (not A300)  and  (not A268) );
 a36340a <=( (not A302)  and  (not A301) );
 a36341a <=( a36340a  and  a36337a );
 a36342a <=( a36341a  and  a36334a );
 a36346a <=( (not A166)  and  (not A167) );
 a36347a <=( (not A169)  and  a36346a );
 a36350a <=( A232  and  A202 );
 a36353a <=( (not A234)  and  A233 );
 a36354a <=( a36353a  and  a36350a );
 a36355a <=( a36354a  and  a36347a );
 a36359a <=( (not A266)  and  (not A265) );
 a36360a <=( (not A235)  and  a36359a );
 a36363a <=( (not A298)  and  (not A268) );
 a36366a <=( (not A301)  and  (not A299) );
 a36367a <=( a36366a  and  a36363a );
 a36368a <=( a36367a  and  a36360a );
 a36372a <=( (not A166)  and  (not A167) );
 a36373a <=( (not A169)  and  a36372a );
 a36376a <=( (not A232)  and  A202 );
 a36379a <=( (not A235)  and  (not A233) );
 a36380a <=( a36379a  and  a36376a );
 a36381a <=( a36380a  and  a36373a );
 a36385a <=( (not A269)  and  (not A268) );
 a36386a <=( (not A267)  and  a36385a );
 a36389a <=( A299  and  A298 );
 a36392a <=( (not A301)  and  (not A300) );
 a36393a <=( a36392a  and  a36389a );
 a36394a <=( a36393a  and  a36386a );
 a36398a <=( (not A166)  and  (not A167) );
 a36399a <=( (not A169)  and  a36398a );
 a36402a <=( (not A232)  and  A202 );
 a36405a <=( (not A235)  and  (not A233) );
 a36406a <=( a36405a  and  a36402a );
 a36407a <=( a36406a  and  a36399a );
 a36411a <=( (not A267)  and  A266 );
 a36412a <=( A265  and  a36411a );
 a36415a <=( (not A300)  and  (not A268) );
 a36418a <=( (not A302)  and  (not A301) );
 a36419a <=( a36418a  and  a36415a );
 a36420a <=( a36419a  and  a36412a );
 a36424a <=( (not A166)  and  (not A167) );
 a36425a <=( (not A169)  and  a36424a );
 a36428a <=( (not A232)  and  A202 );
 a36431a <=( (not A235)  and  (not A233) );
 a36432a <=( a36431a  and  a36428a );
 a36433a <=( a36432a  and  a36425a );
 a36437a <=( (not A267)  and  A266 );
 a36438a <=( A265  and  a36437a );
 a36441a <=( (not A298)  and  (not A268) );
 a36444a <=( (not A301)  and  (not A299) );
 a36445a <=( a36444a  and  a36441a );
 a36446a <=( a36445a  and  a36438a );
 a36450a <=( (not A166)  and  (not A167) );
 a36451a <=( (not A169)  and  a36450a );
 a36454a <=( (not A232)  and  A202 );
 a36457a <=( (not A235)  and  (not A233) );
 a36458a <=( a36457a  and  a36454a );
 a36459a <=( a36458a  and  a36451a );
 a36463a <=( (not A268)  and  (not A266) );
 a36464a <=( (not A265)  and  a36463a );
 a36467a <=( A299  and  A298 );
 a36470a <=( (not A301)  and  (not A300) );
 a36471a <=( a36470a  and  a36467a );
 a36472a <=( a36471a  and  a36464a );
 a36476a <=( (not A166)  and  (not A167) );
 a36477a <=( (not A169)  and  a36476a );
 a36480a <=( A201  and  A199 );
 a36483a <=( (not A235)  and  (not A234) );
 a36484a <=( a36483a  and  a36480a );
 a36485a <=( a36484a  and  a36477a );
 a36489a <=( (not A268)  and  (not A267) );
 a36490a <=( (not A236)  and  a36489a );
 a36493a <=( (not A300)  and  (not A269) );
 a36496a <=( (not A302)  and  (not A301) );
 a36497a <=( a36496a  and  a36493a );
 a36498a <=( a36497a  and  a36490a );
 a36502a <=( (not A166)  and  (not A167) );
 a36503a <=( (not A169)  and  a36502a );
 a36506a <=( A201  and  A199 );
 a36509a <=( (not A235)  and  (not A234) );
 a36510a <=( a36509a  and  a36506a );
 a36511a <=( a36510a  and  a36503a );
 a36515a <=( (not A268)  and  (not A267) );
 a36516a <=( (not A236)  and  a36515a );
 a36519a <=( (not A298)  and  (not A269) );
 a36522a <=( (not A301)  and  (not A299) );
 a36523a <=( a36522a  and  a36519a );
 a36524a <=( a36523a  and  a36516a );
 a36528a <=( (not A166)  and  (not A167) );
 a36529a <=( (not A169)  and  a36528a );
 a36532a <=( A201  and  A199 );
 a36535a <=( (not A235)  and  (not A234) );
 a36536a <=( a36535a  and  a36532a );
 a36537a <=( a36536a  and  a36529a );
 a36541a <=( (not A266)  and  (not A265) );
 a36542a <=( (not A236)  and  a36541a );
 a36545a <=( (not A300)  and  (not A268) );
 a36548a <=( (not A302)  and  (not A301) );
 a36549a <=( a36548a  and  a36545a );
 a36550a <=( a36549a  and  a36542a );
 a36554a <=( (not A166)  and  (not A167) );
 a36555a <=( (not A169)  and  a36554a );
 a36558a <=( A201  and  A199 );
 a36561a <=( (not A235)  and  (not A234) );
 a36562a <=( a36561a  and  a36558a );
 a36563a <=( a36562a  and  a36555a );
 a36567a <=( (not A266)  and  (not A265) );
 a36568a <=( (not A236)  and  a36567a );
 a36571a <=( (not A298)  and  (not A268) );
 a36574a <=( (not A301)  and  (not A299) );
 a36575a <=( a36574a  and  a36571a );
 a36576a <=( a36575a  and  a36568a );
 a36580a <=( (not A166)  and  (not A167) );
 a36581a <=( (not A169)  and  a36580a );
 a36584a <=( A201  and  A199 );
 a36587a <=( (not A233)  and  (not A232) );
 a36588a <=( a36587a  and  a36584a );
 a36589a <=( a36588a  and  a36581a );
 a36593a <=( (not A268)  and  (not A267) );
 a36594a <=( (not A235)  and  a36593a );
 a36597a <=( (not A300)  and  (not A269) );
 a36600a <=( (not A302)  and  (not A301) );
 a36601a <=( a36600a  and  a36597a );
 a36602a <=( a36601a  and  a36594a );
 a36606a <=( (not A166)  and  (not A167) );
 a36607a <=( (not A169)  and  a36606a );
 a36610a <=( A201  and  A199 );
 a36613a <=( (not A233)  and  (not A232) );
 a36614a <=( a36613a  and  a36610a );
 a36615a <=( a36614a  and  a36607a );
 a36619a <=( (not A268)  and  (not A267) );
 a36620a <=( (not A235)  and  a36619a );
 a36623a <=( (not A298)  and  (not A269) );
 a36626a <=( (not A301)  and  (not A299) );
 a36627a <=( a36626a  and  a36623a );
 a36628a <=( a36627a  and  a36620a );
 a36632a <=( (not A166)  and  (not A167) );
 a36633a <=( (not A169)  and  a36632a );
 a36636a <=( A201  and  A199 );
 a36639a <=( (not A233)  and  (not A232) );
 a36640a <=( a36639a  and  a36636a );
 a36641a <=( a36640a  and  a36633a );
 a36645a <=( (not A266)  and  (not A265) );
 a36646a <=( (not A235)  and  a36645a );
 a36649a <=( (not A300)  and  (not A268) );
 a36652a <=( (not A302)  and  (not A301) );
 a36653a <=( a36652a  and  a36649a );
 a36654a <=( a36653a  and  a36646a );
 a36658a <=( (not A166)  and  (not A167) );
 a36659a <=( (not A169)  and  a36658a );
 a36662a <=( A201  and  A199 );
 a36665a <=( (not A233)  and  (not A232) );
 a36666a <=( a36665a  and  a36662a );
 a36667a <=( a36666a  and  a36659a );
 a36671a <=( (not A266)  and  (not A265) );
 a36672a <=( (not A235)  and  a36671a );
 a36675a <=( (not A298)  and  (not A268) );
 a36678a <=( (not A301)  and  (not A299) );
 a36679a <=( a36678a  and  a36675a );
 a36680a <=( a36679a  and  a36672a );
 a36684a <=( (not A166)  and  (not A167) );
 a36685a <=( (not A169)  and  a36684a );
 a36688a <=( A201  and  A200 );
 a36691a <=( (not A235)  and  (not A234) );
 a36692a <=( a36691a  and  a36688a );
 a36693a <=( a36692a  and  a36685a );
 a36697a <=( (not A268)  and  (not A267) );
 a36698a <=( (not A236)  and  a36697a );
 a36701a <=( (not A300)  and  (not A269) );
 a36704a <=( (not A302)  and  (not A301) );
 a36705a <=( a36704a  and  a36701a );
 a36706a <=( a36705a  and  a36698a );
 a36710a <=( (not A166)  and  (not A167) );
 a36711a <=( (not A169)  and  a36710a );
 a36714a <=( A201  and  A200 );
 a36717a <=( (not A235)  and  (not A234) );
 a36718a <=( a36717a  and  a36714a );
 a36719a <=( a36718a  and  a36711a );
 a36723a <=( (not A268)  and  (not A267) );
 a36724a <=( (not A236)  and  a36723a );
 a36727a <=( (not A298)  and  (not A269) );
 a36730a <=( (not A301)  and  (not A299) );
 a36731a <=( a36730a  and  a36727a );
 a36732a <=( a36731a  and  a36724a );
 a36736a <=( (not A166)  and  (not A167) );
 a36737a <=( (not A169)  and  a36736a );
 a36740a <=( A201  and  A200 );
 a36743a <=( (not A235)  and  (not A234) );
 a36744a <=( a36743a  and  a36740a );
 a36745a <=( a36744a  and  a36737a );
 a36749a <=( (not A266)  and  (not A265) );
 a36750a <=( (not A236)  and  a36749a );
 a36753a <=( (not A300)  and  (not A268) );
 a36756a <=( (not A302)  and  (not A301) );
 a36757a <=( a36756a  and  a36753a );
 a36758a <=( a36757a  and  a36750a );
 a36762a <=( (not A166)  and  (not A167) );
 a36763a <=( (not A169)  and  a36762a );
 a36766a <=( A201  and  A200 );
 a36769a <=( (not A235)  and  (not A234) );
 a36770a <=( a36769a  and  a36766a );
 a36771a <=( a36770a  and  a36763a );
 a36775a <=( (not A266)  and  (not A265) );
 a36776a <=( (not A236)  and  a36775a );
 a36779a <=( (not A298)  and  (not A268) );
 a36782a <=( (not A301)  and  (not A299) );
 a36783a <=( a36782a  and  a36779a );
 a36784a <=( a36783a  and  a36776a );
 a36788a <=( (not A166)  and  (not A167) );
 a36789a <=( (not A169)  and  a36788a );
 a36792a <=( A201  and  A200 );
 a36795a <=( (not A233)  and  (not A232) );
 a36796a <=( a36795a  and  a36792a );
 a36797a <=( a36796a  and  a36789a );
 a36801a <=( (not A268)  and  (not A267) );
 a36802a <=( (not A235)  and  a36801a );
 a36805a <=( (not A300)  and  (not A269) );
 a36808a <=( (not A302)  and  (not A301) );
 a36809a <=( a36808a  and  a36805a );
 a36810a <=( a36809a  and  a36802a );
 a36814a <=( (not A166)  and  (not A167) );
 a36815a <=( (not A169)  and  a36814a );
 a36818a <=( A201  and  A200 );
 a36821a <=( (not A233)  and  (not A232) );
 a36822a <=( a36821a  and  a36818a );
 a36823a <=( a36822a  and  a36815a );
 a36827a <=( (not A268)  and  (not A267) );
 a36828a <=( (not A235)  and  a36827a );
 a36831a <=( (not A298)  and  (not A269) );
 a36834a <=( (not A301)  and  (not A299) );
 a36835a <=( a36834a  and  a36831a );
 a36836a <=( a36835a  and  a36828a );
 a36840a <=( (not A166)  and  (not A167) );
 a36841a <=( (not A169)  and  a36840a );
 a36844a <=( A201  and  A200 );
 a36847a <=( (not A233)  and  (not A232) );
 a36848a <=( a36847a  and  a36844a );
 a36849a <=( a36848a  and  a36841a );
 a36853a <=( (not A266)  and  (not A265) );
 a36854a <=( (not A235)  and  a36853a );
 a36857a <=( (not A300)  and  (not A268) );
 a36860a <=( (not A302)  and  (not A301) );
 a36861a <=( a36860a  and  a36857a );
 a36862a <=( a36861a  and  a36854a );
 a36866a <=( (not A166)  and  (not A167) );
 a36867a <=( (not A169)  and  a36866a );
 a36870a <=( A201  and  A200 );
 a36873a <=( (not A233)  and  (not A232) );
 a36874a <=( a36873a  and  a36870a );
 a36875a <=( a36874a  and  a36867a );
 a36879a <=( (not A266)  and  (not A265) );
 a36880a <=( (not A235)  and  a36879a );
 a36883a <=( (not A298)  and  (not A268) );
 a36886a <=( (not A301)  and  (not A299) );
 a36887a <=( a36886a  and  a36883a );
 a36888a <=( a36887a  and  a36880a );
 a36892a <=( A167  and  (not A168) );
 a36893a <=( (not A169)  and  a36892a );
 a36896a <=( A202  and  A166 );
 a36899a <=( (not A235)  and  (not A234) );
 a36900a <=( a36899a  and  a36896a );
 a36901a <=( a36900a  and  a36893a );
 a36905a <=( (not A268)  and  (not A267) );
 a36906a <=( (not A236)  and  a36905a );
 a36909a <=( (not A300)  and  (not A269) );
 a36912a <=( (not A302)  and  (not A301) );
 a36913a <=( a36912a  and  a36909a );
 a36914a <=( a36913a  and  a36906a );
 a36918a <=( A167  and  (not A168) );
 a36919a <=( (not A169)  and  a36918a );
 a36922a <=( A202  and  A166 );
 a36925a <=( (not A235)  and  (not A234) );
 a36926a <=( a36925a  and  a36922a );
 a36927a <=( a36926a  and  a36919a );
 a36931a <=( (not A268)  and  (not A267) );
 a36932a <=( (not A236)  and  a36931a );
 a36935a <=( (not A298)  and  (not A269) );
 a36938a <=( (not A301)  and  (not A299) );
 a36939a <=( a36938a  and  a36935a );
 a36940a <=( a36939a  and  a36932a );
 a36944a <=( A167  and  (not A168) );
 a36945a <=( (not A169)  and  a36944a );
 a36948a <=( A202  and  A166 );
 a36951a <=( (not A235)  and  (not A234) );
 a36952a <=( a36951a  and  a36948a );
 a36953a <=( a36952a  and  a36945a );
 a36957a <=( (not A266)  and  (not A265) );
 a36958a <=( (not A236)  and  a36957a );
 a36961a <=( (not A300)  and  (not A268) );
 a36964a <=( (not A302)  and  (not A301) );
 a36965a <=( a36964a  and  a36961a );
 a36966a <=( a36965a  and  a36958a );
 a36970a <=( A167  and  (not A168) );
 a36971a <=( (not A169)  and  a36970a );
 a36974a <=( A202  and  A166 );
 a36977a <=( (not A235)  and  (not A234) );
 a36978a <=( a36977a  and  a36974a );
 a36979a <=( a36978a  and  a36971a );
 a36983a <=( (not A266)  and  (not A265) );
 a36984a <=( (not A236)  and  a36983a );
 a36987a <=( (not A298)  and  (not A268) );
 a36990a <=( (not A301)  and  (not A299) );
 a36991a <=( a36990a  and  a36987a );
 a36992a <=( a36991a  and  a36984a );
 a36996a <=( A167  and  (not A168) );
 a36997a <=( (not A169)  and  a36996a );
 a37000a <=( A202  and  A166 );
 a37003a <=( (not A233)  and  (not A232) );
 a37004a <=( a37003a  and  a37000a );
 a37005a <=( a37004a  and  a36997a );
 a37009a <=( (not A268)  and  (not A267) );
 a37010a <=( (not A235)  and  a37009a );
 a37013a <=( (not A300)  and  (not A269) );
 a37016a <=( (not A302)  and  (not A301) );
 a37017a <=( a37016a  and  a37013a );
 a37018a <=( a37017a  and  a37010a );
 a37022a <=( A167  and  (not A168) );
 a37023a <=( (not A169)  and  a37022a );
 a37026a <=( A202  and  A166 );
 a37029a <=( (not A233)  and  (not A232) );
 a37030a <=( a37029a  and  a37026a );
 a37031a <=( a37030a  and  a37023a );
 a37035a <=( (not A268)  and  (not A267) );
 a37036a <=( (not A235)  and  a37035a );
 a37039a <=( (not A298)  and  (not A269) );
 a37042a <=( (not A301)  and  (not A299) );
 a37043a <=( a37042a  and  a37039a );
 a37044a <=( a37043a  and  a37036a );
 a37048a <=( A167  and  (not A168) );
 a37049a <=( (not A169)  and  a37048a );
 a37052a <=( A202  and  A166 );
 a37055a <=( (not A233)  and  (not A232) );
 a37056a <=( a37055a  and  a37052a );
 a37057a <=( a37056a  and  a37049a );
 a37061a <=( (not A266)  and  (not A265) );
 a37062a <=( (not A235)  and  a37061a );
 a37065a <=( (not A300)  and  (not A268) );
 a37068a <=( (not A302)  and  (not A301) );
 a37069a <=( a37068a  and  a37065a );
 a37070a <=( a37069a  and  a37062a );
 a37074a <=( A167  and  (not A168) );
 a37075a <=( (not A169)  and  a37074a );
 a37078a <=( A202  and  A166 );
 a37081a <=( (not A233)  and  (not A232) );
 a37082a <=( a37081a  and  a37078a );
 a37083a <=( a37082a  and  a37075a );
 a37087a <=( (not A266)  and  (not A265) );
 a37088a <=( (not A235)  and  a37087a );
 a37091a <=( (not A298)  and  (not A268) );
 a37094a <=( (not A301)  and  (not A299) );
 a37095a <=( a37094a  and  a37091a );
 a37096a <=( a37095a  and  a37088a );
 a37100a <=( (not A168)  and  (not A169) );
 a37101a <=( (not A170)  and  a37100a );
 a37104a <=( (not A234)  and  A202 );
 a37107a <=( (not A236)  and  (not A235) );
 a37108a <=( a37107a  and  a37104a );
 a37109a <=( a37108a  and  a37101a );
 a37113a <=( (not A269)  and  (not A268) );
 a37114a <=( (not A267)  and  a37113a );
 a37117a <=( A299  and  A298 );
 a37120a <=( (not A301)  and  (not A300) );
 a37121a <=( a37120a  and  a37117a );
 a37122a <=( a37121a  and  a37114a );
 a37126a <=( (not A168)  and  (not A169) );
 a37127a <=( (not A170)  and  a37126a );
 a37130a <=( (not A234)  and  A202 );
 a37133a <=( (not A236)  and  (not A235) );
 a37134a <=( a37133a  and  a37130a );
 a37135a <=( a37134a  and  a37127a );
 a37139a <=( (not A267)  and  A266 );
 a37140a <=( A265  and  a37139a );
 a37143a <=( (not A300)  and  (not A268) );
 a37146a <=( (not A302)  and  (not A301) );
 a37147a <=( a37146a  and  a37143a );
 a37148a <=( a37147a  and  a37140a );
 a37152a <=( (not A168)  and  (not A169) );
 a37153a <=( (not A170)  and  a37152a );
 a37156a <=( (not A234)  and  A202 );
 a37159a <=( (not A236)  and  (not A235) );
 a37160a <=( a37159a  and  a37156a );
 a37161a <=( a37160a  and  a37153a );
 a37165a <=( (not A267)  and  A266 );
 a37166a <=( A265  and  a37165a );
 a37169a <=( (not A298)  and  (not A268) );
 a37172a <=( (not A301)  and  (not A299) );
 a37173a <=( a37172a  and  a37169a );
 a37174a <=( a37173a  and  a37166a );
 a37178a <=( (not A168)  and  (not A169) );
 a37179a <=( (not A170)  and  a37178a );
 a37182a <=( (not A234)  and  A202 );
 a37185a <=( (not A236)  and  (not A235) );
 a37186a <=( a37185a  and  a37182a );
 a37187a <=( a37186a  and  a37179a );
 a37191a <=( (not A268)  and  (not A266) );
 a37192a <=( (not A265)  and  a37191a );
 a37195a <=( A299  and  A298 );
 a37198a <=( (not A301)  and  (not A300) );
 a37199a <=( a37198a  and  a37195a );
 a37200a <=( a37199a  and  a37192a );
 a37204a <=( (not A168)  and  (not A169) );
 a37205a <=( (not A170)  and  a37204a );
 a37208a <=( A232  and  A202 );
 a37211a <=( (not A234)  and  A233 );
 a37212a <=( a37211a  and  a37208a );
 a37213a <=( a37212a  and  a37205a );
 a37217a <=( (not A268)  and  (not A267) );
 a37218a <=( (not A235)  and  a37217a );
 a37221a <=( (not A300)  and  (not A269) );
 a37224a <=( (not A302)  and  (not A301) );
 a37225a <=( a37224a  and  a37221a );
 a37226a <=( a37225a  and  a37218a );
 a37230a <=( (not A168)  and  (not A169) );
 a37231a <=( (not A170)  and  a37230a );
 a37234a <=( A232  and  A202 );
 a37237a <=( (not A234)  and  A233 );
 a37238a <=( a37237a  and  a37234a );
 a37239a <=( a37238a  and  a37231a );
 a37243a <=( (not A268)  and  (not A267) );
 a37244a <=( (not A235)  and  a37243a );
 a37247a <=( (not A298)  and  (not A269) );
 a37250a <=( (not A301)  and  (not A299) );
 a37251a <=( a37250a  and  a37247a );
 a37252a <=( a37251a  and  a37244a );
 a37256a <=( (not A168)  and  (not A169) );
 a37257a <=( (not A170)  and  a37256a );
 a37260a <=( A232  and  A202 );
 a37263a <=( (not A234)  and  A233 );
 a37264a <=( a37263a  and  a37260a );
 a37265a <=( a37264a  and  a37257a );
 a37269a <=( (not A266)  and  (not A265) );
 a37270a <=( (not A235)  and  a37269a );
 a37273a <=( (not A300)  and  (not A268) );
 a37276a <=( (not A302)  and  (not A301) );
 a37277a <=( a37276a  and  a37273a );
 a37278a <=( a37277a  and  a37270a );
 a37282a <=( (not A168)  and  (not A169) );
 a37283a <=( (not A170)  and  a37282a );
 a37286a <=( A232  and  A202 );
 a37289a <=( (not A234)  and  A233 );
 a37290a <=( a37289a  and  a37286a );
 a37291a <=( a37290a  and  a37283a );
 a37295a <=( (not A266)  and  (not A265) );
 a37296a <=( (not A235)  and  a37295a );
 a37299a <=( (not A298)  and  (not A268) );
 a37302a <=( (not A301)  and  (not A299) );
 a37303a <=( a37302a  and  a37299a );
 a37304a <=( a37303a  and  a37296a );
 a37308a <=( (not A168)  and  (not A169) );
 a37309a <=( (not A170)  and  a37308a );
 a37312a <=( (not A232)  and  A202 );
 a37315a <=( (not A235)  and  (not A233) );
 a37316a <=( a37315a  and  a37312a );
 a37317a <=( a37316a  and  a37309a );
 a37321a <=( (not A269)  and  (not A268) );
 a37322a <=( (not A267)  and  a37321a );
 a37325a <=( A299  and  A298 );
 a37328a <=( (not A301)  and  (not A300) );
 a37329a <=( a37328a  and  a37325a );
 a37330a <=( a37329a  and  a37322a );
 a37334a <=( (not A168)  and  (not A169) );
 a37335a <=( (not A170)  and  a37334a );
 a37338a <=( (not A232)  and  A202 );
 a37341a <=( (not A235)  and  (not A233) );
 a37342a <=( a37341a  and  a37338a );
 a37343a <=( a37342a  and  a37335a );
 a37347a <=( (not A267)  and  A266 );
 a37348a <=( A265  and  a37347a );
 a37351a <=( (not A300)  and  (not A268) );
 a37354a <=( (not A302)  and  (not A301) );
 a37355a <=( a37354a  and  a37351a );
 a37356a <=( a37355a  and  a37348a );
 a37360a <=( (not A168)  and  (not A169) );
 a37361a <=( (not A170)  and  a37360a );
 a37364a <=( (not A232)  and  A202 );
 a37367a <=( (not A235)  and  (not A233) );
 a37368a <=( a37367a  and  a37364a );
 a37369a <=( a37368a  and  a37361a );
 a37373a <=( (not A267)  and  A266 );
 a37374a <=( A265  and  a37373a );
 a37377a <=( (not A298)  and  (not A268) );
 a37380a <=( (not A301)  and  (not A299) );
 a37381a <=( a37380a  and  a37377a );
 a37382a <=( a37381a  and  a37374a );
 a37386a <=( (not A168)  and  (not A169) );
 a37387a <=( (not A170)  and  a37386a );
 a37390a <=( (not A232)  and  A202 );
 a37393a <=( (not A235)  and  (not A233) );
 a37394a <=( a37393a  and  a37390a );
 a37395a <=( a37394a  and  a37387a );
 a37399a <=( (not A268)  and  (not A266) );
 a37400a <=( (not A265)  and  a37399a );
 a37403a <=( A299  and  A298 );
 a37406a <=( (not A301)  and  (not A300) );
 a37407a <=( a37406a  and  a37403a );
 a37408a <=( a37407a  and  a37400a );
 a37412a <=( (not A168)  and  (not A169) );
 a37413a <=( (not A170)  and  a37412a );
 a37416a <=( A201  and  A199 );
 a37419a <=( (not A235)  and  (not A234) );
 a37420a <=( a37419a  and  a37416a );
 a37421a <=( a37420a  and  a37413a );
 a37425a <=( (not A268)  and  (not A267) );
 a37426a <=( (not A236)  and  a37425a );
 a37429a <=( (not A300)  and  (not A269) );
 a37432a <=( (not A302)  and  (not A301) );
 a37433a <=( a37432a  and  a37429a );
 a37434a <=( a37433a  and  a37426a );
 a37438a <=( (not A168)  and  (not A169) );
 a37439a <=( (not A170)  and  a37438a );
 a37442a <=( A201  and  A199 );
 a37445a <=( (not A235)  and  (not A234) );
 a37446a <=( a37445a  and  a37442a );
 a37447a <=( a37446a  and  a37439a );
 a37451a <=( (not A268)  and  (not A267) );
 a37452a <=( (not A236)  and  a37451a );
 a37455a <=( (not A298)  and  (not A269) );
 a37458a <=( (not A301)  and  (not A299) );
 a37459a <=( a37458a  and  a37455a );
 a37460a <=( a37459a  and  a37452a );
 a37464a <=( (not A168)  and  (not A169) );
 a37465a <=( (not A170)  and  a37464a );
 a37468a <=( A201  and  A199 );
 a37471a <=( (not A235)  and  (not A234) );
 a37472a <=( a37471a  and  a37468a );
 a37473a <=( a37472a  and  a37465a );
 a37477a <=( (not A266)  and  (not A265) );
 a37478a <=( (not A236)  and  a37477a );
 a37481a <=( (not A300)  and  (not A268) );
 a37484a <=( (not A302)  and  (not A301) );
 a37485a <=( a37484a  and  a37481a );
 a37486a <=( a37485a  and  a37478a );
 a37490a <=( (not A168)  and  (not A169) );
 a37491a <=( (not A170)  and  a37490a );
 a37494a <=( A201  and  A199 );
 a37497a <=( (not A235)  and  (not A234) );
 a37498a <=( a37497a  and  a37494a );
 a37499a <=( a37498a  and  a37491a );
 a37503a <=( (not A266)  and  (not A265) );
 a37504a <=( (not A236)  and  a37503a );
 a37507a <=( (not A298)  and  (not A268) );
 a37510a <=( (not A301)  and  (not A299) );
 a37511a <=( a37510a  and  a37507a );
 a37512a <=( a37511a  and  a37504a );
 a37516a <=( (not A168)  and  (not A169) );
 a37517a <=( (not A170)  and  a37516a );
 a37520a <=( A201  and  A199 );
 a37523a <=( (not A233)  and  (not A232) );
 a37524a <=( a37523a  and  a37520a );
 a37525a <=( a37524a  and  a37517a );
 a37529a <=( (not A268)  and  (not A267) );
 a37530a <=( (not A235)  and  a37529a );
 a37533a <=( (not A300)  and  (not A269) );
 a37536a <=( (not A302)  and  (not A301) );
 a37537a <=( a37536a  and  a37533a );
 a37538a <=( a37537a  and  a37530a );
 a37542a <=( (not A168)  and  (not A169) );
 a37543a <=( (not A170)  and  a37542a );
 a37546a <=( A201  and  A199 );
 a37549a <=( (not A233)  and  (not A232) );
 a37550a <=( a37549a  and  a37546a );
 a37551a <=( a37550a  and  a37543a );
 a37555a <=( (not A268)  and  (not A267) );
 a37556a <=( (not A235)  and  a37555a );
 a37559a <=( (not A298)  and  (not A269) );
 a37562a <=( (not A301)  and  (not A299) );
 a37563a <=( a37562a  and  a37559a );
 a37564a <=( a37563a  and  a37556a );
 a37568a <=( (not A168)  and  (not A169) );
 a37569a <=( (not A170)  and  a37568a );
 a37572a <=( A201  and  A199 );
 a37575a <=( (not A233)  and  (not A232) );
 a37576a <=( a37575a  and  a37572a );
 a37577a <=( a37576a  and  a37569a );
 a37581a <=( (not A266)  and  (not A265) );
 a37582a <=( (not A235)  and  a37581a );
 a37585a <=( (not A300)  and  (not A268) );
 a37588a <=( (not A302)  and  (not A301) );
 a37589a <=( a37588a  and  a37585a );
 a37590a <=( a37589a  and  a37582a );
 a37594a <=( (not A168)  and  (not A169) );
 a37595a <=( (not A170)  and  a37594a );
 a37598a <=( A201  and  A199 );
 a37601a <=( (not A233)  and  (not A232) );
 a37602a <=( a37601a  and  a37598a );
 a37603a <=( a37602a  and  a37595a );
 a37607a <=( (not A266)  and  (not A265) );
 a37608a <=( (not A235)  and  a37607a );
 a37611a <=( (not A298)  and  (not A268) );
 a37614a <=( (not A301)  and  (not A299) );
 a37615a <=( a37614a  and  a37611a );
 a37616a <=( a37615a  and  a37608a );
 a37620a <=( (not A168)  and  (not A169) );
 a37621a <=( (not A170)  and  a37620a );
 a37624a <=( A201  and  A200 );
 a37627a <=( (not A235)  and  (not A234) );
 a37628a <=( a37627a  and  a37624a );
 a37629a <=( a37628a  and  a37621a );
 a37633a <=( (not A268)  and  (not A267) );
 a37634a <=( (not A236)  and  a37633a );
 a37637a <=( (not A300)  and  (not A269) );
 a37640a <=( (not A302)  and  (not A301) );
 a37641a <=( a37640a  and  a37637a );
 a37642a <=( a37641a  and  a37634a );
 a37646a <=( (not A168)  and  (not A169) );
 a37647a <=( (not A170)  and  a37646a );
 a37650a <=( A201  and  A200 );
 a37653a <=( (not A235)  and  (not A234) );
 a37654a <=( a37653a  and  a37650a );
 a37655a <=( a37654a  and  a37647a );
 a37659a <=( (not A268)  and  (not A267) );
 a37660a <=( (not A236)  and  a37659a );
 a37663a <=( (not A298)  and  (not A269) );
 a37666a <=( (not A301)  and  (not A299) );
 a37667a <=( a37666a  and  a37663a );
 a37668a <=( a37667a  and  a37660a );
 a37672a <=( (not A168)  and  (not A169) );
 a37673a <=( (not A170)  and  a37672a );
 a37676a <=( A201  and  A200 );
 a37679a <=( (not A235)  and  (not A234) );
 a37680a <=( a37679a  and  a37676a );
 a37681a <=( a37680a  and  a37673a );
 a37685a <=( (not A266)  and  (not A265) );
 a37686a <=( (not A236)  and  a37685a );
 a37689a <=( (not A300)  and  (not A268) );
 a37692a <=( (not A302)  and  (not A301) );
 a37693a <=( a37692a  and  a37689a );
 a37694a <=( a37693a  and  a37686a );
 a37698a <=( (not A168)  and  (not A169) );
 a37699a <=( (not A170)  and  a37698a );
 a37702a <=( A201  and  A200 );
 a37705a <=( (not A235)  and  (not A234) );
 a37706a <=( a37705a  and  a37702a );
 a37707a <=( a37706a  and  a37699a );
 a37711a <=( (not A266)  and  (not A265) );
 a37712a <=( (not A236)  and  a37711a );
 a37715a <=( (not A298)  and  (not A268) );
 a37718a <=( (not A301)  and  (not A299) );
 a37719a <=( a37718a  and  a37715a );
 a37720a <=( a37719a  and  a37712a );
 a37724a <=( (not A168)  and  (not A169) );
 a37725a <=( (not A170)  and  a37724a );
 a37728a <=( A201  and  A200 );
 a37731a <=( (not A233)  and  (not A232) );
 a37732a <=( a37731a  and  a37728a );
 a37733a <=( a37732a  and  a37725a );
 a37737a <=( (not A268)  and  (not A267) );
 a37738a <=( (not A235)  and  a37737a );
 a37741a <=( (not A300)  and  (not A269) );
 a37744a <=( (not A302)  and  (not A301) );
 a37745a <=( a37744a  and  a37741a );
 a37746a <=( a37745a  and  a37738a );
 a37750a <=( (not A168)  and  (not A169) );
 a37751a <=( (not A170)  and  a37750a );
 a37754a <=( A201  and  A200 );
 a37757a <=( (not A233)  and  (not A232) );
 a37758a <=( a37757a  and  a37754a );
 a37759a <=( a37758a  and  a37751a );
 a37763a <=( (not A268)  and  (not A267) );
 a37764a <=( (not A235)  and  a37763a );
 a37767a <=( (not A298)  and  (not A269) );
 a37770a <=( (not A301)  and  (not A299) );
 a37771a <=( a37770a  and  a37767a );
 a37772a <=( a37771a  and  a37764a );
 a37776a <=( (not A168)  and  (not A169) );
 a37777a <=( (not A170)  and  a37776a );
 a37780a <=( A201  and  A200 );
 a37783a <=( (not A233)  and  (not A232) );
 a37784a <=( a37783a  and  a37780a );
 a37785a <=( a37784a  and  a37777a );
 a37789a <=( (not A266)  and  (not A265) );
 a37790a <=( (not A235)  and  a37789a );
 a37793a <=( (not A300)  and  (not A268) );
 a37796a <=( (not A302)  and  (not A301) );
 a37797a <=( a37796a  and  a37793a );
 a37798a <=( a37797a  and  a37790a );
 a37802a <=( (not A168)  and  (not A169) );
 a37803a <=( (not A170)  and  a37802a );
 a37806a <=( A201  and  A200 );
 a37809a <=( (not A233)  and  (not A232) );
 a37810a <=( a37809a  and  a37806a );
 a37811a <=( a37810a  and  a37803a );
 a37815a <=( (not A266)  and  (not A265) );
 a37816a <=( (not A235)  and  a37815a );
 a37819a <=( (not A298)  and  (not A268) );
 a37822a <=( (not A301)  and  (not A299) );
 a37823a <=( a37822a  and  a37819a );
 a37824a <=( a37823a  and  a37816a );
 a37828a <=( (not A201)  and  A166 );
 a37829a <=( A168  and  a37828a );
 a37832a <=( (not A203)  and  (not A202) );
 a37835a <=( (not A235)  and  (not A234) );
 a37836a <=( a37835a  and  a37832a );
 a37837a <=( a37836a  and  a37829a );
 a37840a <=( (not A267)  and  (not A236) );
 a37843a <=( (not A269)  and  (not A268) );
 a37844a <=( a37843a  and  a37840a );
 a37847a <=( A299  and  A298 );
 a37850a <=( (not A301)  and  (not A300) );
 a37851a <=( a37850a  and  a37847a );
 a37852a <=( a37851a  and  a37844a );
 a37856a <=( (not A201)  and  A166 );
 a37857a <=( A168  and  a37856a );
 a37860a <=( (not A203)  and  (not A202) );
 a37863a <=( (not A235)  and  (not A234) );
 a37864a <=( a37863a  and  a37860a );
 a37865a <=( a37864a  and  a37857a );
 a37868a <=( A265  and  (not A236) );
 a37871a <=( (not A267)  and  A266 );
 a37872a <=( a37871a  and  a37868a );
 a37875a <=( (not A300)  and  (not A268) );
 a37878a <=( (not A302)  and  (not A301) );
 a37879a <=( a37878a  and  a37875a );
 a37880a <=( a37879a  and  a37872a );
 a37884a <=( (not A201)  and  A166 );
 a37885a <=( A168  and  a37884a );
 a37888a <=( (not A203)  and  (not A202) );
 a37891a <=( (not A235)  and  (not A234) );
 a37892a <=( a37891a  and  a37888a );
 a37893a <=( a37892a  and  a37885a );
 a37896a <=( A265  and  (not A236) );
 a37899a <=( (not A267)  and  A266 );
 a37900a <=( a37899a  and  a37896a );
 a37903a <=( (not A298)  and  (not A268) );
 a37906a <=( (not A301)  and  (not A299) );
 a37907a <=( a37906a  and  a37903a );
 a37908a <=( a37907a  and  a37900a );
 a37912a <=( (not A201)  and  A166 );
 a37913a <=( A168  and  a37912a );
 a37916a <=( (not A203)  and  (not A202) );
 a37919a <=( (not A235)  and  (not A234) );
 a37920a <=( a37919a  and  a37916a );
 a37921a <=( a37920a  and  a37913a );
 a37924a <=( (not A265)  and  (not A236) );
 a37927a <=( (not A268)  and  (not A266) );
 a37928a <=( a37927a  and  a37924a );
 a37931a <=( A299  and  A298 );
 a37934a <=( (not A301)  and  (not A300) );
 a37935a <=( a37934a  and  a37931a );
 a37936a <=( a37935a  and  a37928a );
 a37940a <=( (not A201)  and  A166 );
 a37941a <=( A168  and  a37940a );
 a37944a <=( (not A203)  and  (not A202) );
 a37947a <=( A233  and  A232 );
 a37948a <=( a37947a  and  a37944a );
 a37949a <=( a37948a  and  a37941a );
 a37952a <=( (not A235)  and  (not A234) );
 a37955a <=( (not A268)  and  (not A267) );
 a37956a <=( a37955a  and  a37952a );
 a37959a <=( (not A300)  and  (not A269) );
 a37962a <=( (not A302)  and  (not A301) );
 a37963a <=( a37962a  and  a37959a );
 a37964a <=( a37963a  and  a37956a );
 a37968a <=( (not A201)  and  A166 );
 a37969a <=( A168  and  a37968a );
 a37972a <=( (not A203)  and  (not A202) );
 a37975a <=( A233  and  A232 );
 a37976a <=( a37975a  and  a37972a );
 a37977a <=( a37976a  and  a37969a );
 a37980a <=( (not A235)  and  (not A234) );
 a37983a <=( (not A268)  and  (not A267) );
 a37984a <=( a37983a  and  a37980a );
 a37987a <=( (not A298)  and  (not A269) );
 a37990a <=( (not A301)  and  (not A299) );
 a37991a <=( a37990a  and  a37987a );
 a37992a <=( a37991a  and  a37984a );
 a37996a <=( (not A201)  and  A166 );
 a37997a <=( A168  and  a37996a );
 a38000a <=( (not A203)  and  (not A202) );
 a38003a <=( A233  and  A232 );
 a38004a <=( a38003a  and  a38000a );
 a38005a <=( a38004a  and  a37997a );
 a38008a <=( (not A235)  and  (not A234) );
 a38011a <=( (not A266)  and  (not A265) );
 a38012a <=( a38011a  and  a38008a );
 a38015a <=( (not A300)  and  (not A268) );
 a38018a <=( (not A302)  and  (not A301) );
 a38019a <=( a38018a  and  a38015a );
 a38020a <=( a38019a  and  a38012a );
 a38024a <=( (not A201)  and  A166 );
 a38025a <=( A168  and  a38024a );
 a38028a <=( (not A203)  and  (not A202) );
 a38031a <=( A233  and  A232 );
 a38032a <=( a38031a  and  a38028a );
 a38033a <=( a38032a  and  a38025a );
 a38036a <=( (not A235)  and  (not A234) );
 a38039a <=( (not A266)  and  (not A265) );
 a38040a <=( a38039a  and  a38036a );
 a38043a <=( (not A298)  and  (not A268) );
 a38046a <=( (not A301)  and  (not A299) );
 a38047a <=( a38046a  and  a38043a );
 a38048a <=( a38047a  and  a38040a );
 a38052a <=( (not A201)  and  A166 );
 a38053a <=( A168  and  a38052a );
 a38056a <=( (not A203)  and  (not A202) );
 a38059a <=( (not A233)  and  (not A232) );
 a38060a <=( a38059a  and  a38056a );
 a38061a <=( a38060a  and  a38053a );
 a38064a <=( (not A267)  and  (not A235) );
 a38067a <=( (not A269)  and  (not A268) );
 a38068a <=( a38067a  and  a38064a );
 a38071a <=( A299  and  A298 );
 a38074a <=( (not A301)  and  (not A300) );
 a38075a <=( a38074a  and  a38071a );
 a38076a <=( a38075a  and  a38068a );
 a38080a <=( (not A201)  and  A166 );
 a38081a <=( A168  and  a38080a );
 a38084a <=( (not A203)  and  (not A202) );
 a38087a <=( (not A233)  and  (not A232) );
 a38088a <=( a38087a  and  a38084a );
 a38089a <=( a38088a  and  a38081a );
 a38092a <=( A265  and  (not A235) );
 a38095a <=( (not A267)  and  A266 );
 a38096a <=( a38095a  and  a38092a );
 a38099a <=( (not A300)  and  (not A268) );
 a38102a <=( (not A302)  and  (not A301) );
 a38103a <=( a38102a  and  a38099a );
 a38104a <=( a38103a  and  a38096a );
 a38108a <=( (not A201)  and  A166 );
 a38109a <=( A168  and  a38108a );
 a38112a <=( (not A203)  and  (not A202) );
 a38115a <=( (not A233)  and  (not A232) );
 a38116a <=( a38115a  and  a38112a );
 a38117a <=( a38116a  and  a38109a );
 a38120a <=( A265  and  (not A235) );
 a38123a <=( (not A267)  and  A266 );
 a38124a <=( a38123a  and  a38120a );
 a38127a <=( (not A298)  and  (not A268) );
 a38130a <=( (not A301)  and  (not A299) );
 a38131a <=( a38130a  and  a38127a );
 a38132a <=( a38131a  and  a38124a );
 a38136a <=( (not A201)  and  A166 );
 a38137a <=( A168  and  a38136a );
 a38140a <=( (not A203)  and  (not A202) );
 a38143a <=( (not A233)  and  (not A232) );
 a38144a <=( a38143a  and  a38140a );
 a38145a <=( a38144a  and  a38137a );
 a38148a <=( (not A265)  and  (not A235) );
 a38151a <=( (not A268)  and  (not A266) );
 a38152a <=( a38151a  and  a38148a );
 a38155a <=( A299  and  A298 );
 a38158a <=( (not A301)  and  (not A300) );
 a38159a <=( a38158a  and  a38155a );
 a38160a <=( a38159a  and  a38152a );
 a38164a <=( A199  and  A166 );
 a38165a <=( A168  and  a38164a );
 a38168a <=( (not A201)  and  A200 );
 a38171a <=( (not A234)  and  (not A202) );
 a38172a <=( a38171a  and  a38168a );
 a38173a <=( a38172a  and  a38165a );
 a38176a <=( (not A236)  and  (not A235) );
 a38179a <=( (not A268)  and  (not A267) );
 a38180a <=( a38179a  and  a38176a );
 a38183a <=( (not A300)  and  (not A269) );
 a38186a <=( (not A302)  and  (not A301) );
 a38187a <=( a38186a  and  a38183a );
 a38188a <=( a38187a  and  a38180a );
 a38192a <=( A199  and  A166 );
 a38193a <=( A168  and  a38192a );
 a38196a <=( (not A201)  and  A200 );
 a38199a <=( (not A234)  and  (not A202) );
 a38200a <=( a38199a  and  a38196a );
 a38201a <=( a38200a  and  a38193a );
 a38204a <=( (not A236)  and  (not A235) );
 a38207a <=( (not A268)  and  (not A267) );
 a38208a <=( a38207a  and  a38204a );
 a38211a <=( (not A298)  and  (not A269) );
 a38214a <=( (not A301)  and  (not A299) );
 a38215a <=( a38214a  and  a38211a );
 a38216a <=( a38215a  and  a38208a );
 a38220a <=( A199  and  A166 );
 a38221a <=( A168  and  a38220a );
 a38224a <=( (not A201)  and  A200 );
 a38227a <=( (not A234)  and  (not A202) );
 a38228a <=( a38227a  and  a38224a );
 a38229a <=( a38228a  and  a38221a );
 a38232a <=( (not A236)  and  (not A235) );
 a38235a <=( (not A266)  and  (not A265) );
 a38236a <=( a38235a  and  a38232a );
 a38239a <=( (not A300)  and  (not A268) );
 a38242a <=( (not A302)  and  (not A301) );
 a38243a <=( a38242a  and  a38239a );
 a38244a <=( a38243a  and  a38236a );
 a38248a <=( A199  and  A166 );
 a38249a <=( A168  and  a38248a );
 a38252a <=( (not A201)  and  A200 );
 a38255a <=( (not A234)  and  (not A202) );
 a38256a <=( a38255a  and  a38252a );
 a38257a <=( a38256a  and  a38249a );
 a38260a <=( (not A236)  and  (not A235) );
 a38263a <=( (not A266)  and  (not A265) );
 a38264a <=( a38263a  and  a38260a );
 a38267a <=( (not A298)  and  (not A268) );
 a38270a <=( (not A301)  and  (not A299) );
 a38271a <=( a38270a  and  a38267a );
 a38272a <=( a38271a  and  a38264a );
 a38276a <=( A199  and  A166 );
 a38277a <=( A168  and  a38276a );
 a38280a <=( (not A201)  and  A200 );
 a38283a <=( (not A232)  and  (not A202) );
 a38284a <=( a38283a  and  a38280a );
 a38285a <=( a38284a  and  a38277a );
 a38288a <=( (not A235)  and  (not A233) );
 a38291a <=( (not A268)  and  (not A267) );
 a38292a <=( a38291a  and  a38288a );
 a38295a <=( (not A300)  and  (not A269) );
 a38298a <=( (not A302)  and  (not A301) );
 a38299a <=( a38298a  and  a38295a );
 a38300a <=( a38299a  and  a38292a );
 a38304a <=( A199  and  A166 );
 a38305a <=( A168  and  a38304a );
 a38308a <=( (not A201)  and  A200 );
 a38311a <=( (not A232)  and  (not A202) );
 a38312a <=( a38311a  and  a38308a );
 a38313a <=( a38312a  and  a38305a );
 a38316a <=( (not A235)  and  (not A233) );
 a38319a <=( (not A268)  and  (not A267) );
 a38320a <=( a38319a  and  a38316a );
 a38323a <=( (not A298)  and  (not A269) );
 a38326a <=( (not A301)  and  (not A299) );
 a38327a <=( a38326a  and  a38323a );
 a38328a <=( a38327a  and  a38320a );
 a38332a <=( A199  and  A166 );
 a38333a <=( A168  and  a38332a );
 a38336a <=( (not A201)  and  A200 );
 a38339a <=( (not A232)  and  (not A202) );
 a38340a <=( a38339a  and  a38336a );
 a38341a <=( a38340a  and  a38333a );
 a38344a <=( (not A235)  and  (not A233) );
 a38347a <=( (not A266)  and  (not A265) );
 a38348a <=( a38347a  and  a38344a );
 a38351a <=( (not A300)  and  (not A268) );
 a38354a <=( (not A302)  and  (not A301) );
 a38355a <=( a38354a  and  a38351a );
 a38356a <=( a38355a  and  a38348a );
 a38360a <=( A199  and  A166 );
 a38361a <=( A168  and  a38360a );
 a38364a <=( (not A201)  and  A200 );
 a38367a <=( (not A232)  and  (not A202) );
 a38368a <=( a38367a  and  a38364a );
 a38369a <=( a38368a  and  a38361a );
 a38372a <=( (not A235)  and  (not A233) );
 a38375a <=( (not A266)  and  (not A265) );
 a38376a <=( a38375a  and  a38372a );
 a38379a <=( (not A298)  and  (not A268) );
 a38382a <=( (not A301)  and  (not A299) );
 a38383a <=( a38382a  and  a38379a );
 a38384a <=( a38383a  and  a38376a );
 a38388a <=( (not A199)  and  A166 );
 a38389a <=( A168  and  a38388a );
 a38392a <=( (not A202)  and  (not A200) );
 a38395a <=( (not A235)  and  (not A234) );
 a38396a <=( a38395a  and  a38392a );
 a38397a <=( a38396a  and  a38389a );
 a38400a <=( (not A267)  and  (not A236) );
 a38403a <=( (not A269)  and  (not A268) );
 a38404a <=( a38403a  and  a38400a );
 a38407a <=( A299  and  A298 );
 a38410a <=( (not A301)  and  (not A300) );
 a38411a <=( a38410a  and  a38407a );
 a38412a <=( a38411a  and  a38404a );
 a38416a <=( (not A199)  and  A166 );
 a38417a <=( A168  and  a38416a );
 a38420a <=( (not A202)  and  (not A200) );
 a38423a <=( (not A235)  and  (not A234) );
 a38424a <=( a38423a  and  a38420a );
 a38425a <=( a38424a  and  a38417a );
 a38428a <=( A265  and  (not A236) );
 a38431a <=( (not A267)  and  A266 );
 a38432a <=( a38431a  and  a38428a );
 a38435a <=( (not A300)  and  (not A268) );
 a38438a <=( (not A302)  and  (not A301) );
 a38439a <=( a38438a  and  a38435a );
 a38440a <=( a38439a  and  a38432a );
 a38444a <=( (not A199)  and  A166 );
 a38445a <=( A168  and  a38444a );
 a38448a <=( (not A202)  and  (not A200) );
 a38451a <=( (not A235)  and  (not A234) );
 a38452a <=( a38451a  and  a38448a );
 a38453a <=( a38452a  and  a38445a );
 a38456a <=( A265  and  (not A236) );
 a38459a <=( (not A267)  and  A266 );
 a38460a <=( a38459a  and  a38456a );
 a38463a <=( (not A298)  and  (not A268) );
 a38466a <=( (not A301)  and  (not A299) );
 a38467a <=( a38466a  and  a38463a );
 a38468a <=( a38467a  and  a38460a );
 a38472a <=( (not A199)  and  A166 );
 a38473a <=( A168  and  a38472a );
 a38476a <=( (not A202)  and  (not A200) );
 a38479a <=( (not A235)  and  (not A234) );
 a38480a <=( a38479a  and  a38476a );
 a38481a <=( a38480a  and  a38473a );
 a38484a <=( (not A265)  and  (not A236) );
 a38487a <=( (not A268)  and  (not A266) );
 a38488a <=( a38487a  and  a38484a );
 a38491a <=( A299  and  A298 );
 a38494a <=( (not A301)  and  (not A300) );
 a38495a <=( a38494a  and  a38491a );
 a38496a <=( a38495a  and  a38488a );
 a38500a <=( (not A199)  and  A166 );
 a38501a <=( A168  and  a38500a );
 a38504a <=( (not A202)  and  (not A200) );
 a38507a <=( A233  and  A232 );
 a38508a <=( a38507a  and  a38504a );
 a38509a <=( a38508a  and  a38501a );
 a38512a <=( (not A235)  and  (not A234) );
 a38515a <=( (not A268)  and  (not A267) );
 a38516a <=( a38515a  and  a38512a );
 a38519a <=( (not A300)  and  (not A269) );
 a38522a <=( (not A302)  and  (not A301) );
 a38523a <=( a38522a  and  a38519a );
 a38524a <=( a38523a  and  a38516a );
 a38528a <=( (not A199)  and  A166 );
 a38529a <=( A168  and  a38528a );
 a38532a <=( (not A202)  and  (not A200) );
 a38535a <=( A233  and  A232 );
 a38536a <=( a38535a  and  a38532a );
 a38537a <=( a38536a  and  a38529a );
 a38540a <=( (not A235)  and  (not A234) );
 a38543a <=( (not A268)  and  (not A267) );
 a38544a <=( a38543a  and  a38540a );
 a38547a <=( (not A298)  and  (not A269) );
 a38550a <=( (not A301)  and  (not A299) );
 a38551a <=( a38550a  and  a38547a );
 a38552a <=( a38551a  and  a38544a );
 a38556a <=( (not A199)  and  A166 );
 a38557a <=( A168  and  a38556a );
 a38560a <=( (not A202)  and  (not A200) );
 a38563a <=( A233  and  A232 );
 a38564a <=( a38563a  and  a38560a );
 a38565a <=( a38564a  and  a38557a );
 a38568a <=( (not A235)  and  (not A234) );
 a38571a <=( (not A266)  and  (not A265) );
 a38572a <=( a38571a  and  a38568a );
 a38575a <=( (not A300)  and  (not A268) );
 a38578a <=( (not A302)  and  (not A301) );
 a38579a <=( a38578a  and  a38575a );
 a38580a <=( a38579a  and  a38572a );
 a38584a <=( (not A199)  and  A166 );
 a38585a <=( A168  and  a38584a );
 a38588a <=( (not A202)  and  (not A200) );
 a38591a <=( A233  and  A232 );
 a38592a <=( a38591a  and  a38588a );
 a38593a <=( a38592a  and  a38585a );
 a38596a <=( (not A235)  and  (not A234) );
 a38599a <=( (not A266)  and  (not A265) );
 a38600a <=( a38599a  and  a38596a );
 a38603a <=( (not A298)  and  (not A268) );
 a38606a <=( (not A301)  and  (not A299) );
 a38607a <=( a38606a  and  a38603a );
 a38608a <=( a38607a  and  a38600a );
 a38612a <=( (not A199)  and  A166 );
 a38613a <=( A168  and  a38612a );
 a38616a <=( (not A202)  and  (not A200) );
 a38619a <=( (not A233)  and  (not A232) );
 a38620a <=( a38619a  and  a38616a );
 a38621a <=( a38620a  and  a38613a );
 a38624a <=( (not A267)  and  (not A235) );
 a38627a <=( (not A269)  and  (not A268) );
 a38628a <=( a38627a  and  a38624a );
 a38631a <=( A299  and  A298 );
 a38634a <=( (not A301)  and  (not A300) );
 a38635a <=( a38634a  and  a38631a );
 a38636a <=( a38635a  and  a38628a );
 a38640a <=( (not A199)  and  A166 );
 a38641a <=( A168  and  a38640a );
 a38644a <=( (not A202)  and  (not A200) );
 a38647a <=( (not A233)  and  (not A232) );
 a38648a <=( a38647a  and  a38644a );
 a38649a <=( a38648a  and  a38641a );
 a38652a <=( A265  and  (not A235) );
 a38655a <=( (not A267)  and  A266 );
 a38656a <=( a38655a  and  a38652a );
 a38659a <=( (not A300)  and  (not A268) );
 a38662a <=( (not A302)  and  (not A301) );
 a38663a <=( a38662a  and  a38659a );
 a38664a <=( a38663a  and  a38656a );
 a38668a <=( (not A199)  and  A166 );
 a38669a <=( A168  and  a38668a );
 a38672a <=( (not A202)  and  (not A200) );
 a38675a <=( (not A233)  and  (not A232) );
 a38676a <=( a38675a  and  a38672a );
 a38677a <=( a38676a  and  a38669a );
 a38680a <=( A265  and  (not A235) );
 a38683a <=( (not A267)  and  A266 );
 a38684a <=( a38683a  and  a38680a );
 a38687a <=( (not A298)  and  (not A268) );
 a38690a <=( (not A301)  and  (not A299) );
 a38691a <=( a38690a  and  a38687a );
 a38692a <=( a38691a  and  a38684a );
 a38696a <=( (not A199)  and  A166 );
 a38697a <=( A168  and  a38696a );
 a38700a <=( (not A202)  and  (not A200) );
 a38703a <=( (not A233)  and  (not A232) );
 a38704a <=( a38703a  and  a38700a );
 a38705a <=( a38704a  and  a38697a );
 a38708a <=( (not A265)  and  (not A235) );
 a38711a <=( (not A268)  and  (not A266) );
 a38712a <=( a38711a  and  a38708a );
 a38715a <=( A299  and  A298 );
 a38718a <=( (not A301)  and  (not A300) );
 a38719a <=( a38718a  and  a38715a );
 a38720a <=( a38719a  and  a38712a );
 a38724a <=( (not A201)  and  A167 );
 a38725a <=( A168  and  a38724a );
 a38728a <=( (not A203)  and  (not A202) );
 a38731a <=( (not A235)  and  (not A234) );
 a38732a <=( a38731a  and  a38728a );
 a38733a <=( a38732a  and  a38725a );
 a38736a <=( (not A267)  and  (not A236) );
 a38739a <=( (not A269)  and  (not A268) );
 a38740a <=( a38739a  and  a38736a );
 a38743a <=( A299  and  A298 );
 a38746a <=( (not A301)  and  (not A300) );
 a38747a <=( a38746a  and  a38743a );
 a38748a <=( a38747a  and  a38740a );
 a38752a <=( (not A201)  and  A167 );
 a38753a <=( A168  and  a38752a );
 a38756a <=( (not A203)  and  (not A202) );
 a38759a <=( (not A235)  and  (not A234) );
 a38760a <=( a38759a  and  a38756a );
 a38761a <=( a38760a  and  a38753a );
 a38764a <=( A265  and  (not A236) );
 a38767a <=( (not A267)  and  A266 );
 a38768a <=( a38767a  and  a38764a );
 a38771a <=( (not A300)  and  (not A268) );
 a38774a <=( (not A302)  and  (not A301) );
 a38775a <=( a38774a  and  a38771a );
 a38776a <=( a38775a  and  a38768a );
 a38780a <=( (not A201)  and  A167 );
 a38781a <=( A168  and  a38780a );
 a38784a <=( (not A203)  and  (not A202) );
 a38787a <=( (not A235)  and  (not A234) );
 a38788a <=( a38787a  and  a38784a );
 a38789a <=( a38788a  and  a38781a );
 a38792a <=( A265  and  (not A236) );
 a38795a <=( (not A267)  and  A266 );
 a38796a <=( a38795a  and  a38792a );
 a38799a <=( (not A298)  and  (not A268) );
 a38802a <=( (not A301)  and  (not A299) );
 a38803a <=( a38802a  and  a38799a );
 a38804a <=( a38803a  and  a38796a );
 a38808a <=( (not A201)  and  A167 );
 a38809a <=( A168  and  a38808a );
 a38812a <=( (not A203)  and  (not A202) );
 a38815a <=( (not A235)  and  (not A234) );
 a38816a <=( a38815a  and  a38812a );
 a38817a <=( a38816a  and  a38809a );
 a38820a <=( (not A265)  and  (not A236) );
 a38823a <=( (not A268)  and  (not A266) );
 a38824a <=( a38823a  and  a38820a );
 a38827a <=( A299  and  A298 );
 a38830a <=( (not A301)  and  (not A300) );
 a38831a <=( a38830a  and  a38827a );
 a38832a <=( a38831a  and  a38824a );
 a38836a <=( (not A201)  and  A167 );
 a38837a <=( A168  and  a38836a );
 a38840a <=( (not A203)  and  (not A202) );
 a38843a <=( A233  and  A232 );
 a38844a <=( a38843a  and  a38840a );
 a38845a <=( a38844a  and  a38837a );
 a38848a <=( (not A235)  and  (not A234) );
 a38851a <=( (not A268)  and  (not A267) );
 a38852a <=( a38851a  and  a38848a );
 a38855a <=( (not A300)  and  (not A269) );
 a38858a <=( (not A302)  and  (not A301) );
 a38859a <=( a38858a  and  a38855a );
 a38860a <=( a38859a  and  a38852a );
 a38864a <=( (not A201)  and  A167 );
 a38865a <=( A168  and  a38864a );
 a38868a <=( (not A203)  and  (not A202) );
 a38871a <=( A233  and  A232 );
 a38872a <=( a38871a  and  a38868a );
 a38873a <=( a38872a  and  a38865a );
 a38876a <=( (not A235)  and  (not A234) );
 a38879a <=( (not A268)  and  (not A267) );
 a38880a <=( a38879a  and  a38876a );
 a38883a <=( (not A298)  and  (not A269) );
 a38886a <=( (not A301)  and  (not A299) );
 a38887a <=( a38886a  and  a38883a );
 a38888a <=( a38887a  and  a38880a );
 a38892a <=( (not A201)  and  A167 );
 a38893a <=( A168  and  a38892a );
 a38896a <=( (not A203)  and  (not A202) );
 a38899a <=( A233  and  A232 );
 a38900a <=( a38899a  and  a38896a );
 a38901a <=( a38900a  and  a38893a );
 a38904a <=( (not A235)  and  (not A234) );
 a38907a <=( (not A266)  and  (not A265) );
 a38908a <=( a38907a  and  a38904a );
 a38911a <=( (not A300)  and  (not A268) );
 a38914a <=( (not A302)  and  (not A301) );
 a38915a <=( a38914a  and  a38911a );
 a38916a <=( a38915a  and  a38908a );
 a38920a <=( (not A201)  and  A167 );
 a38921a <=( A168  and  a38920a );
 a38924a <=( (not A203)  and  (not A202) );
 a38927a <=( A233  and  A232 );
 a38928a <=( a38927a  and  a38924a );
 a38929a <=( a38928a  and  a38921a );
 a38932a <=( (not A235)  and  (not A234) );
 a38935a <=( (not A266)  and  (not A265) );
 a38936a <=( a38935a  and  a38932a );
 a38939a <=( (not A298)  and  (not A268) );
 a38942a <=( (not A301)  and  (not A299) );
 a38943a <=( a38942a  and  a38939a );
 a38944a <=( a38943a  and  a38936a );
 a38948a <=( (not A201)  and  A167 );
 a38949a <=( A168  and  a38948a );
 a38952a <=( (not A203)  and  (not A202) );
 a38955a <=( (not A233)  and  (not A232) );
 a38956a <=( a38955a  and  a38952a );
 a38957a <=( a38956a  and  a38949a );
 a38960a <=( (not A267)  and  (not A235) );
 a38963a <=( (not A269)  and  (not A268) );
 a38964a <=( a38963a  and  a38960a );
 a38967a <=( A299  and  A298 );
 a38970a <=( (not A301)  and  (not A300) );
 a38971a <=( a38970a  and  a38967a );
 a38972a <=( a38971a  and  a38964a );
 a38976a <=( (not A201)  and  A167 );
 a38977a <=( A168  and  a38976a );
 a38980a <=( (not A203)  and  (not A202) );
 a38983a <=( (not A233)  and  (not A232) );
 a38984a <=( a38983a  and  a38980a );
 a38985a <=( a38984a  and  a38977a );
 a38988a <=( A265  and  (not A235) );
 a38991a <=( (not A267)  and  A266 );
 a38992a <=( a38991a  and  a38988a );
 a38995a <=( (not A300)  and  (not A268) );
 a38998a <=( (not A302)  and  (not A301) );
 a38999a <=( a38998a  and  a38995a );
 a39000a <=( a38999a  and  a38992a );
 a39004a <=( (not A201)  and  A167 );
 a39005a <=( A168  and  a39004a );
 a39008a <=( (not A203)  and  (not A202) );
 a39011a <=( (not A233)  and  (not A232) );
 a39012a <=( a39011a  and  a39008a );
 a39013a <=( a39012a  and  a39005a );
 a39016a <=( A265  and  (not A235) );
 a39019a <=( (not A267)  and  A266 );
 a39020a <=( a39019a  and  a39016a );
 a39023a <=( (not A298)  and  (not A268) );
 a39026a <=( (not A301)  and  (not A299) );
 a39027a <=( a39026a  and  a39023a );
 a39028a <=( a39027a  and  a39020a );
 a39032a <=( (not A201)  and  A167 );
 a39033a <=( A168  and  a39032a );
 a39036a <=( (not A203)  and  (not A202) );
 a39039a <=( (not A233)  and  (not A232) );
 a39040a <=( a39039a  and  a39036a );
 a39041a <=( a39040a  and  a39033a );
 a39044a <=( (not A265)  and  (not A235) );
 a39047a <=( (not A268)  and  (not A266) );
 a39048a <=( a39047a  and  a39044a );
 a39051a <=( A299  and  A298 );
 a39054a <=( (not A301)  and  (not A300) );
 a39055a <=( a39054a  and  a39051a );
 a39056a <=( a39055a  and  a39048a );
 a39060a <=( A199  and  A167 );
 a39061a <=( A168  and  a39060a );
 a39064a <=( (not A201)  and  A200 );
 a39067a <=( (not A234)  and  (not A202) );
 a39068a <=( a39067a  and  a39064a );
 a39069a <=( a39068a  and  a39061a );
 a39072a <=( (not A236)  and  (not A235) );
 a39075a <=( (not A268)  and  (not A267) );
 a39076a <=( a39075a  and  a39072a );
 a39079a <=( (not A300)  and  (not A269) );
 a39082a <=( (not A302)  and  (not A301) );
 a39083a <=( a39082a  and  a39079a );
 a39084a <=( a39083a  and  a39076a );
 a39088a <=( A199  and  A167 );
 a39089a <=( A168  and  a39088a );
 a39092a <=( (not A201)  and  A200 );
 a39095a <=( (not A234)  and  (not A202) );
 a39096a <=( a39095a  and  a39092a );
 a39097a <=( a39096a  and  a39089a );
 a39100a <=( (not A236)  and  (not A235) );
 a39103a <=( (not A268)  and  (not A267) );
 a39104a <=( a39103a  and  a39100a );
 a39107a <=( (not A298)  and  (not A269) );
 a39110a <=( (not A301)  and  (not A299) );
 a39111a <=( a39110a  and  a39107a );
 a39112a <=( a39111a  and  a39104a );
 a39116a <=( A199  and  A167 );
 a39117a <=( A168  and  a39116a );
 a39120a <=( (not A201)  and  A200 );
 a39123a <=( (not A234)  and  (not A202) );
 a39124a <=( a39123a  and  a39120a );
 a39125a <=( a39124a  and  a39117a );
 a39128a <=( (not A236)  and  (not A235) );
 a39131a <=( (not A266)  and  (not A265) );
 a39132a <=( a39131a  and  a39128a );
 a39135a <=( (not A300)  and  (not A268) );
 a39138a <=( (not A302)  and  (not A301) );
 a39139a <=( a39138a  and  a39135a );
 a39140a <=( a39139a  and  a39132a );
 a39144a <=( A199  and  A167 );
 a39145a <=( A168  and  a39144a );
 a39148a <=( (not A201)  and  A200 );
 a39151a <=( (not A234)  and  (not A202) );
 a39152a <=( a39151a  and  a39148a );
 a39153a <=( a39152a  and  a39145a );
 a39156a <=( (not A236)  and  (not A235) );
 a39159a <=( (not A266)  and  (not A265) );
 a39160a <=( a39159a  and  a39156a );
 a39163a <=( (not A298)  and  (not A268) );
 a39166a <=( (not A301)  and  (not A299) );
 a39167a <=( a39166a  and  a39163a );
 a39168a <=( a39167a  and  a39160a );
 a39172a <=( A199  and  A167 );
 a39173a <=( A168  and  a39172a );
 a39176a <=( (not A201)  and  A200 );
 a39179a <=( (not A232)  and  (not A202) );
 a39180a <=( a39179a  and  a39176a );
 a39181a <=( a39180a  and  a39173a );
 a39184a <=( (not A235)  and  (not A233) );
 a39187a <=( (not A268)  and  (not A267) );
 a39188a <=( a39187a  and  a39184a );
 a39191a <=( (not A300)  and  (not A269) );
 a39194a <=( (not A302)  and  (not A301) );
 a39195a <=( a39194a  and  a39191a );
 a39196a <=( a39195a  and  a39188a );
 a39200a <=( A199  and  A167 );
 a39201a <=( A168  and  a39200a );
 a39204a <=( (not A201)  and  A200 );
 a39207a <=( (not A232)  and  (not A202) );
 a39208a <=( a39207a  and  a39204a );
 a39209a <=( a39208a  and  a39201a );
 a39212a <=( (not A235)  and  (not A233) );
 a39215a <=( (not A268)  and  (not A267) );
 a39216a <=( a39215a  and  a39212a );
 a39219a <=( (not A298)  and  (not A269) );
 a39222a <=( (not A301)  and  (not A299) );
 a39223a <=( a39222a  and  a39219a );
 a39224a <=( a39223a  and  a39216a );
 a39228a <=( A199  and  A167 );
 a39229a <=( A168  and  a39228a );
 a39232a <=( (not A201)  and  A200 );
 a39235a <=( (not A232)  and  (not A202) );
 a39236a <=( a39235a  and  a39232a );
 a39237a <=( a39236a  and  a39229a );
 a39240a <=( (not A235)  and  (not A233) );
 a39243a <=( (not A266)  and  (not A265) );
 a39244a <=( a39243a  and  a39240a );
 a39247a <=( (not A300)  and  (not A268) );
 a39250a <=( (not A302)  and  (not A301) );
 a39251a <=( a39250a  and  a39247a );
 a39252a <=( a39251a  and  a39244a );
 a39256a <=( A199  and  A167 );
 a39257a <=( A168  and  a39256a );
 a39260a <=( (not A201)  and  A200 );
 a39263a <=( (not A232)  and  (not A202) );
 a39264a <=( a39263a  and  a39260a );
 a39265a <=( a39264a  and  a39257a );
 a39268a <=( (not A235)  and  (not A233) );
 a39271a <=( (not A266)  and  (not A265) );
 a39272a <=( a39271a  and  a39268a );
 a39275a <=( (not A298)  and  (not A268) );
 a39278a <=( (not A301)  and  (not A299) );
 a39279a <=( a39278a  and  a39275a );
 a39280a <=( a39279a  and  a39272a );
 a39284a <=( (not A199)  and  A167 );
 a39285a <=( A168  and  a39284a );
 a39288a <=( (not A202)  and  (not A200) );
 a39291a <=( (not A235)  and  (not A234) );
 a39292a <=( a39291a  and  a39288a );
 a39293a <=( a39292a  and  a39285a );
 a39296a <=( (not A267)  and  (not A236) );
 a39299a <=( (not A269)  and  (not A268) );
 a39300a <=( a39299a  and  a39296a );
 a39303a <=( A299  and  A298 );
 a39306a <=( (not A301)  and  (not A300) );
 a39307a <=( a39306a  and  a39303a );
 a39308a <=( a39307a  and  a39300a );
 a39312a <=( (not A199)  and  A167 );
 a39313a <=( A168  and  a39312a );
 a39316a <=( (not A202)  and  (not A200) );
 a39319a <=( (not A235)  and  (not A234) );
 a39320a <=( a39319a  and  a39316a );
 a39321a <=( a39320a  and  a39313a );
 a39324a <=( A265  and  (not A236) );
 a39327a <=( (not A267)  and  A266 );
 a39328a <=( a39327a  and  a39324a );
 a39331a <=( (not A300)  and  (not A268) );
 a39334a <=( (not A302)  and  (not A301) );
 a39335a <=( a39334a  and  a39331a );
 a39336a <=( a39335a  and  a39328a );
 a39340a <=( (not A199)  and  A167 );
 a39341a <=( A168  and  a39340a );
 a39344a <=( (not A202)  and  (not A200) );
 a39347a <=( (not A235)  and  (not A234) );
 a39348a <=( a39347a  and  a39344a );
 a39349a <=( a39348a  and  a39341a );
 a39352a <=( A265  and  (not A236) );
 a39355a <=( (not A267)  and  A266 );
 a39356a <=( a39355a  and  a39352a );
 a39359a <=( (not A298)  and  (not A268) );
 a39362a <=( (not A301)  and  (not A299) );
 a39363a <=( a39362a  and  a39359a );
 a39364a <=( a39363a  and  a39356a );
 a39368a <=( (not A199)  and  A167 );
 a39369a <=( A168  and  a39368a );
 a39372a <=( (not A202)  and  (not A200) );
 a39375a <=( (not A235)  and  (not A234) );
 a39376a <=( a39375a  and  a39372a );
 a39377a <=( a39376a  and  a39369a );
 a39380a <=( (not A265)  and  (not A236) );
 a39383a <=( (not A268)  and  (not A266) );
 a39384a <=( a39383a  and  a39380a );
 a39387a <=( A299  and  A298 );
 a39390a <=( (not A301)  and  (not A300) );
 a39391a <=( a39390a  and  a39387a );
 a39392a <=( a39391a  and  a39384a );
 a39396a <=( (not A199)  and  A167 );
 a39397a <=( A168  and  a39396a );
 a39400a <=( (not A202)  and  (not A200) );
 a39403a <=( A233  and  A232 );
 a39404a <=( a39403a  and  a39400a );
 a39405a <=( a39404a  and  a39397a );
 a39408a <=( (not A235)  and  (not A234) );
 a39411a <=( (not A268)  and  (not A267) );
 a39412a <=( a39411a  and  a39408a );
 a39415a <=( (not A300)  and  (not A269) );
 a39418a <=( (not A302)  and  (not A301) );
 a39419a <=( a39418a  and  a39415a );
 a39420a <=( a39419a  and  a39412a );
 a39424a <=( (not A199)  and  A167 );
 a39425a <=( A168  and  a39424a );
 a39428a <=( (not A202)  and  (not A200) );
 a39431a <=( A233  and  A232 );
 a39432a <=( a39431a  and  a39428a );
 a39433a <=( a39432a  and  a39425a );
 a39436a <=( (not A235)  and  (not A234) );
 a39439a <=( (not A268)  and  (not A267) );
 a39440a <=( a39439a  and  a39436a );
 a39443a <=( (not A298)  and  (not A269) );
 a39446a <=( (not A301)  and  (not A299) );
 a39447a <=( a39446a  and  a39443a );
 a39448a <=( a39447a  and  a39440a );
 a39452a <=( (not A199)  and  A167 );
 a39453a <=( A168  and  a39452a );
 a39456a <=( (not A202)  and  (not A200) );
 a39459a <=( A233  and  A232 );
 a39460a <=( a39459a  and  a39456a );
 a39461a <=( a39460a  and  a39453a );
 a39464a <=( (not A235)  and  (not A234) );
 a39467a <=( (not A266)  and  (not A265) );
 a39468a <=( a39467a  and  a39464a );
 a39471a <=( (not A300)  and  (not A268) );
 a39474a <=( (not A302)  and  (not A301) );
 a39475a <=( a39474a  and  a39471a );
 a39476a <=( a39475a  and  a39468a );
 a39480a <=( (not A199)  and  A167 );
 a39481a <=( A168  and  a39480a );
 a39484a <=( (not A202)  and  (not A200) );
 a39487a <=( A233  and  A232 );
 a39488a <=( a39487a  and  a39484a );
 a39489a <=( a39488a  and  a39481a );
 a39492a <=( (not A235)  and  (not A234) );
 a39495a <=( (not A266)  and  (not A265) );
 a39496a <=( a39495a  and  a39492a );
 a39499a <=( (not A298)  and  (not A268) );
 a39502a <=( (not A301)  and  (not A299) );
 a39503a <=( a39502a  and  a39499a );
 a39504a <=( a39503a  and  a39496a );
 a39508a <=( (not A199)  and  A167 );
 a39509a <=( A168  and  a39508a );
 a39512a <=( (not A202)  and  (not A200) );
 a39515a <=( (not A233)  and  (not A232) );
 a39516a <=( a39515a  and  a39512a );
 a39517a <=( a39516a  and  a39509a );
 a39520a <=( (not A267)  and  (not A235) );
 a39523a <=( (not A269)  and  (not A268) );
 a39524a <=( a39523a  and  a39520a );
 a39527a <=( A299  and  A298 );
 a39530a <=( (not A301)  and  (not A300) );
 a39531a <=( a39530a  and  a39527a );
 a39532a <=( a39531a  and  a39524a );
 a39536a <=( (not A199)  and  A167 );
 a39537a <=( A168  and  a39536a );
 a39540a <=( (not A202)  and  (not A200) );
 a39543a <=( (not A233)  and  (not A232) );
 a39544a <=( a39543a  and  a39540a );
 a39545a <=( a39544a  and  a39537a );
 a39548a <=( A265  and  (not A235) );
 a39551a <=( (not A267)  and  A266 );
 a39552a <=( a39551a  and  a39548a );
 a39555a <=( (not A300)  and  (not A268) );
 a39558a <=( (not A302)  and  (not A301) );
 a39559a <=( a39558a  and  a39555a );
 a39560a <=( a39559a  and  a39552a );
 a39564a <=( (not A199)  and  A167 );
 a39565a <=( A168  and  a39564a );
 a39568a <=( (not A202)  and  (not A200) );
 a39571a <=( (not A233)  and  (not A232) );
 a39572a <=( a39571a  and  a39568a );
 a39573a <=( a39572a  and  a39565a );
 a39576a <=( A265  and  (not A235) );
 a39579a <=( (not A267)  and  A266 );
 a39580a <=( a39579a  and  a39576a );
 a39583a <=( (not A298)  and  (not A268) );
 a39586a <=( (not A301)  and  (not A299) );
 a39587a <=( a39586a  and  a39583a );
 a39588a <=( a39587a  and  a39580a );
 a39592a <=( (not A199)  and  A167 );
 a39593a <=( A168  and  a39592a );
 a39596a <=( (not A202)  and  (not A200) );
 a39599a <=( (not A233)  and  (not A232) );
 a39600a <=( a39599a  and  a39596a );
 a39601a <=( a39600a  and  a39593a );
 a39604a <=( (not A265)  and  (not A235) );
 a39607a <=( (not A268)  and  (not A266) );
 a39608a <=( a39607a  and  a39604a );
 a39611a <=( A299  and  A298 );
 a39614a <=( (not A301)  and  (not A300) );
 a39615a <=( a39614a  and  a39611a );
 a39616a <=( a39615a  and  a39608a );
 a39620a <=( (not A166)  and  A167 );
 a39621a <=( A170  and  a39620a );
 a39624a <=( (not A202)  and  (not A201) );
 a39627a <=( (not A234)  and  (not A203) );
 a39628a <=( a39627a  and  a39624a );
 a39629a <=( a39628a  and  a39621a );
 a39632a <=( (not A236)  and  (not A235) );
 a39635a <=( (not A268)  and  (not A267) );
 a39636a <=( a39635a  and  a39632a );
 a39639a <=( (not A300)  and  (not A269) );
 a39642a <=( (not A302)  and  (not A301) );
 a39643a <=( a39642a  and  a39639a );
 a39644a <=( a39643a  and  a39636a );
 a39648a <=( (not A166)  and  A167 );
 a39649a <=( A170  and  a39648a );
 a39652a <=( (not A202)  and  (not A201) );
 a39655a <=( (not A234)  and  (not A203) );
 a39656a <=( a39655a  and  a39652a );
 a39657a <=( a39656a  and  a39649a );
 a39660a <=( (not A236)  and  (not A235) );
 a39663a <=( (not A268)  and  (not A267) );
 a39664a <=( a39663a  and  a39660a );
 a39667a <=( (not A298)  and  (not A269) );
 a39670a <=( (not A301)  and  (not A299) );
 a39671a <=( a39670a  and  a39667a );
 a39672a <=( a39671a  and  a39664a );
 a39676a <=( (not A166)  and  A167 );
 a39677a <=( A170  and  a39676a );
 a39680a <=( (not A202)  and  (not A201) );
 a39683a <=( (not A234)  and  (not A203) );
 a39684a <=( a39683a  and  a39680a );
 a39685a <=( a39684a  and  a39677a );
 a39688a <=( (not A236)  and  (not A235) );
 a39691a <=( (not A266)  and  (not A265) );
 a39692a <=( a39691a  and  a39688a );
 a39695a <=( (not A300)  and  (not A268) );
 a39698a <=( (not A302)  and  (not A301) );
 a39699a <=( a39698a  and  a39695a );
 a39700a <=( a39699a  and  a39692a );
 a39704a <=( (not A166)  and  A167 );
 a39705a <=( A170  and  a39704a );
 a39708a <=( (not A202)  and  (not A201) );
 a39711a <=( (not A234)  and  (not A203) );
 a39712a <=( a39711a  and  a39708a );
 a39713a <=( a39712a  and  a39705a );
 a39716a <=( (not A236)  and  (not A235) );
 a39719a <=( (not A266)  and  (not A265) );
 a39720a <=( a39719a  and  a39716a );
 a39723a <=( (not A298)  and  (not A268) );
 a39726a <=( (not A301)  and  (not A299) );
 a39727a <=( a39726a  and  a39723a );
 a39728a <=( a39727a  and  a39720a );
 a39732a <=( (not A166)  and  A167 );
 a39733a <=( A170  and  a39732a );
 a39736a <=( (not A202)  and  (not A201) );
 a39739a <=( (not A232)  and  (not A203) );
 a39740a <=( a39739a  and  a39736a );
 a39741a <=( a39740a  and  a39733a );
 a39744a <=( (not A235)  and  (not A233) );
 a39747a <=( (not A268)  and  (not A267) );
 a39748a <=( a39747a  and  a39744a );
 a39751a <=( (not A300)  and  (not A269) );
 a39754a <=( (not A302)  and  (not A301) );
 a39755a <=( a39754a  and  a39751a );
 a39756a <=( a39755a  and  a39748a );
 a39760a <=( (not A166)  and  A167 );
 a39761a <=( A170  and  a39760a );
 a39764a <=( (not A202)  and  (not A201) );
 a39767a <=( (not A232)  and  (not A203) );
 a39768a <=( a39767a  and  a39764a );
 a39769a <=( a39768a  and  a39761a );
 a39772a <=( (not A235)  and  (not A233) );
 a39775a <=( (not A268)  and  (not A267) );
 a39776a <=( a39775a  and  a39772a );
 a39779a <=( (not A298)  and  (not A269) );
 a39782a <=( (not A301)  and  (not A299) );
 a39783a <=( a39782a  and  a39779a );
 a39784a <=( a39783a  and  a39776a );
 a39788a <=( (not A166)  and  A167 );
 a39789a <=( A170  and  a39788a );
 a39792a <=( (not A202)  and  (not A201) );
 a39795a <=( (not A232)  and  (not A203) );
 a39796a <=( a39795a  and  a39792a );
 a39797a <=( a39796a  and  a39789a );
 a39800a <=( (not A235)  and  (not A233) );
 a39803a <=( (not A266)  and  (not A265) );
 a39804a <=( a39803a  and  a39800a );
 a39807a <=( (not A300)  and  (not A268) );
 a39810a <=( (not A302)  and  (not A301) );
 a39811a <=( a39810a  and  a39807a );
 a39812a <=( a39811a  and  a39804a );
 a39816a <=( (not A166)  and  A167 );
 a39817a <=( A170  and  a39816a );
 a39820a <=( (not A202)  and  (not A201) );
 a39823a <=( (not A232)  and  (not A203) );
 a39824a <=( a39823a  and  a39820a );
 a39825a <=( a39824a  and  a39817a );
 a39828a <=( (not A235)  and  (not A233) );
 a39831a <=( (not A266)  and  (not A265) );
 a39832a <=( a39831a  and  a39828a );
 a39835a <=( (not A298)  and  (not A268) );
 a39838a <=( (not A301)  and  (not A299) );
 a39839a <=( a39838a  and  a39835a );
 a39840a <=( a39839a  and  a39832a );
 a39844a <=( (not A166)  and  A167 );
 a39845a <=( A170  and  a39844a );
 a39848a <=( (not A200)  and  (not A199) );
 a39851a <=( (not A234)  and  (not A202) );
 a39852a <=( a39851a  and  a39848a );
 a39853a <=( a39852a  and  a39845a );
 a39856a <=( (not A236)  and  (not A235) );
 a39859a <=( (not A268)  and  (not A267) );
 a39860a <=( a39859a  and  a39856a );
 a39863a <=( (not A300)  and  (not A269) );
 a39866a <=( (not A302)  and  (not A301) );
 a39867a <=( a39866a  and  a39863a );
 a39868a <=( a39867a  and  a39860a );
 a39872a <=( (not A166)  and  A167 );
 a39873a <=( A170  and  a39872a );
 a39876a <=( (not A200)  and  (not A199) );
 a39879a <=( (not A234)  and  (not A202) );
 a39880a <=( a39879a  and  a39876a );
 a39881a <=( a39880a  and  a39873a );
 a39884a <=( (not A236)  and  (not A235) );
 a39887a <=( (not A268)  and  (not A267) );
 a39888a <=( a39887a  and  a39884a );
 a39891a <=( (not A298)  and  (not A269) );
 a39894a <=( (not A301)  and  (not A299) );
 a39895a <=( a39894a  and  a39891a );
 a39896a <=( a39895a  and  a39888a );
 a39900a <=( (not A166)  and  A167 );
 a39901a <=( A170  and  a39900a );
 a39904a <=( (not A200)  and  (not A199) );
 a39907a <=( (not A234)  and  (not A202) );
 a39908a <=( a39907a  and  a39904a );
 a39909a <=( a39908a  and  a39901a );
 a39912a <=( (not A236)  and  (not A235) );
 a39915a <=( (not A266)  and  (not A265) );
 a39916a <=( a39915a  and  a39912a );
 a39919a <=( (not A300)  and  (not A268) );
 a39922a <=( (not A302)  and  (not A301) );
 a39923a <=( a39922a  and  a39919a );
 a39924a <=( a39923a  and  a39916a );
 a39928a <=( (not A166)  and  A167 );
 a39929a <=( A170  and  a39928a );
 a39932a <=( (not A200)  and  (not A199) );
 a39935a <=( (not A234)  and  (not A202) );
 a39936a <=( a39935a  and  a39932a );
 a39937a <=( a39936a  and  a39929a );
 a39940a <=( (not A236)  and  (not A235) );
 a39943a <=( (not A266)  and  (not A265) );
 a39944a <=( a39943a  and  a39940a );
 a39947a <=( (not A298)  and  (not A268) );
 a39950a <=( (not A301)  and  (not A299) );
 a39951a <=( a39950a  and  a39947a );
 a39952a <=( a39951a  and  a39944a );
 a39956a <=( (not A166)  and  A167 );
 a39957a <=( A170  and  a39956a );
 a39960a <=( (not A200)  and  (not A199) );
 a39963a <=( (not A232)  and  (not A202) );
 a39964a <=( a39963a  and  a39960a );
 a39965a <=( a39964a  and  a39957a );
 a39968a <=( (not A235)  and  (not A233) );
 a39971a <=( (not A268)  and  (not A267) );
 a39972a <=( a39971a  and  a39968a );
 a39975a <=( (not A300)  and  (not A269) );
 a39978a <=( (not A302)  and  (not A301) );
 a39979a <=( a39978a  and  a39975a );
 a39980a <=( a39979a  and  a39972a );
 a39984a <=( (not A166)  and  A167 );
 a39985a <=( A170  and  a39984a );
 a39988a <=( (not A200)  and  (not A199) );
 a39991a <=( (not A232)  and  (not A202) );
 a39992a <=( a39991a  and  a39988a );
 a39993a <=( a39992a  and  a39985a );
 a39996a <=( (not A235)  and  (not A233) );
 a39999a <=( (not A268)  and  (not A267) );
 a40000a <=( a39999a  and  a39996a );
 a40003a <=( (not A298)  and  (not A269) );
 a40006a <=( (not A301)  and  (not A299) );
 a40007a <=( a40006a  and  a40003a );
 a40008a <=( a40007a  and  a40000a );
 a40012a <=( (not A166)  and  A167 );
 a40013a <=( A170  and  a40012a );
 a40016a <=( (not A200)  and  (not A199) );
 a40019a <=( (not A232)  and  (not A202) );
 a40020a <=( a40019a  and  a40016a );
 a40021a <=( a40020a  and  a40013a );
 a40024a <=( (not A235)  and  (not A233) );
 a40027a <=( (not A266)  and  (not A265) );
 a40028a <=( a40027a  and  a40024a );
 a40031a <=( (not A300)  and  (not A268) );
 a40034a <=( (not A302)  and  (not A301) );
 a40035a <=( a40034a  and  a40031a );
 a40036a <=( a40035a  and  a40028a );
 a40040a <=( (not A166)  and  A167 );
 a40041a <=( A170  and  a40040a );
 a40044a <=( (not A200)  and  (not A199) );
 a40047a <=( (not A232)  and  (not A202) );
 a40048a <=( a40047a  and  a40044a );
 a40049a <=( a40048a  and  a40041a );
 a40052a <=( (not A235)  and  (not A233) );
 a40055a <=( (not A266)  and  (not A265) );
 a40056a <=( a40055a  and  a40052a );
 a40059a <=( (not A298)  and  (not A268) );
 a40062a <=( (not A301)  and  (not A299) );
 a40063a <=( a40062a  and  a40059a );
 a40064a <=( a40063a  and  a40056a );
 a40068a <=( A166  and  (not A167) );
 a40069a <=( A170  and  a40068a );
 a40072a <=( (not A202)  and  (not A201) );
 a40075a <=( (not A234)  and  (not A203) );
 a40076a <=( a40075a  and  a40072a );
 a40077a <=( a40076a  and  a40069a );
 a40080a <=( (not A236)  and  (not A235) );
 a40083a <=( (not A268)  and  (not A267) );
 a40084a <=( a40083a  and  a40080a );
 a40087a <=( (not A300)  and  (not A269) );
 a40090a <=( (not A302)  and  (not A301) );
 a40091a <=( a40090a  and  a40087a );
 a40092a <=( a40091a  and  a40084a );
 a40096a <=( A166  and  (not A167) );
 a40097a <=( A170  and  a40096a );
 a40100a <=( (not A202)  and  (not A201) );
 a40103a <=( (not A234)  and  (not A203) );
 a40104a <=( a40103a  and  a40100a );
 a40105a <=( a40104a  and  a40097a );
 a40108a <=( (not A236)  and  (not A235) );
 a40111a <=( (not A268)  and  (not A267) );
 a40112a <=( a40111a  and  a40108a );
 a40115a <=( (not A298)  and  (not A269) );
 a40118a <=( (not A301)  and  (not A299) );
 a40119a <=( a40118a  and  a40115a );
 a40120a <=( a40119a  and  a40112a );
 a40124a <=( A166  and  (not A167) );
 a40125a <=( A170  and  a40124a );
 a40128a <=( (not A202)  and  (not A201) );
 a40131a <=( (not A234)  and  (not A203) );
 a40132a <=( a40131a  and  a40128a );
 a40133a <=( a40132a  and  a40125a );
 a40136a <=( (not A236)  and  (not A235) );
 a40139a <=( (not A266)  and  (not A265) );
 a40140a <=( a40139a  and  a40136a );
 a40143a <=( (not A300)  and  (not A268) );
 a40146a <=( (not A302)  and  (not A301) );
 a40147a <=( a40146a  and  a40143a );
 a40148a <=( a40147a  and  a40140a );
 a40152a <=( A166  and  (not A167) );
 a40153a <=( A170  and  a40152a );
 a40156a <=( (not A202)  and  (not A201) );
 a40159a <=( (not A234)  and  (not A203) );
 a40160a <=( a40159a  and  a40156a );
 a40161a <=( a40160a  and  a40153a );
 a40164a <=( (not A236)  and  (not A235) );
 a40167a <=( (not A266)  and  (not A265) );
 a40168a <=( a40167a  and  a40164a );
 a40171a <=( (not A298)  and  (not A268) );
 a40174a <=( (not A301)  and  (not A299) );
 a40175a <=( a40174a  and  a40171a );
 a40176a <=( a40175a  and  a40168a );
 a40180a <=( A166  and  (not A167) );
 a40181a <=( A170  and  a40180a );
 a40184a <=( (not A202)  and  (not A201) );
 a40187a <=( (not A232)  and  (not A203) );
 a40188a <=( a40187a  and  a40184a );
 a40189a <=( a40188a  and  a40181a );
 a40192a <=( (not A235)  and  (not A233) );
 a40195a <=( (not A268)  and  (not A267) );
 a40196a <=( a40195a  and  a40192a );
 a40199a <=( (not A300)  and  (not A269) );
 a40202a <=( (not A302)  and  (not A301) );
 a40203a <=( a40202a  and  a40199a );
 a40204a <=( a40203a  and  a40196a );
 a40208a <=( A166  and  (not A167) );
 a40209a <=( A170  and  a40208a );
 a40212a <=( (not A202)  and  (not A201) );
 a40215a <=( (not A232)  and  (not A203) );
 a40216a <=( a40215a  and  a40212a );
 a40217a <=( a40216a  and  a40209a );
 a40220a <=( (not A235)  and  (not A233) );
 a40223a <=( (not A268)  and  (not A267) );
 a40224a <=( a40223a  and  a40220a );
 a40227a <=( (not A298)  and  (not A269) );
 a40230a <=( (not A301)  and  (not A299) );
 a40231a <=( a40230a  and  a40227a );
 a40232a <=( a40231a  and  a40224a );
 a40236a <=( A166  and  (not A167) );
 a40237a <=( A170  and  a40236a );
 a40240a <=( (not A202)  and  (not A201) );
 a40243a <=( (not A232)  and  (not A203) );
 a40244a <=( a40243a  and  a40240a );
 a40245a <=( a40244a  and  a40237a );
 a40248a <=( (not A235)  and  (not A233) );
 a40251a <=( (not A266)  and  (not A265) );
 a40252a <=( a40251a  and  a40248a );
 a40255a <=( (not A300)  and  (not A268) );
 a40258a <=( (not A302)  and  (not A301) );
 a40259a <=( a40258a  and  a40255a );
 a40260a <=( a40259a  and  a40252a );
 a40264a <=( A166  and  (not A167) );
 a40265a <=( A170  and  a40264a );
 a40268a <=( (not A202)  and  (not A201) );
 a40271a <=( (not A232)  and  (not A203) );
 a40272a <=( a40271a  and  a40268a );
 a40273a <=( a40272a  and  a40265a );
 a40276a <=( (not A235)  and  (not A233) );
 a40279a <=( (not A266)  and  (not A265) );
 a40280a <=( a40279a  and  a40276a );
 a40283a <=( (not A298)  and  (not A268) );
 a40286a <=( (not A301)  and  (not A299) );
 a40287a <=( a40286a  and  a40283a );
 a40288a <=( a40287a  and  a40280a );
 a40292a <=( A166  and  (not A167) );
 a40293a <=( A170  and  a40292a );
 a40296a <=( (not A200)  and  (not A199) );
 a40299a <=( (not A234)  and  (not A202) );
 a40300a <=( a40299a  and  a40296a );
 a40301a <=( a40300a  and  a40293a );
 a40304a <=( (not A236)  and  (not A235) );
 a40307a <=( (not A268)  and  (not A267) );
 a40308a <=( a40307a  and  a40304a );
 a40311a <=( (not A300)  and  (not A269) );
 a40314a <=( (not A302)  and  (not A301) );
 a40315a <=( a40314a  and  a40311a );
 a40316a <=( a40315a  and  a40308a );
 a40320a <=( A166  and  (not A167) );
 a40321a <=( A170  and  a40320a );
 a40324a <=( (not A200)  and  (not A199) );
 a40327a <=( (not A234)  and  (not A202) );
 a40328a <=( a40327a  and  a40324a );
 a40329a <=( a40328a  and  a40321a );
 a40332a <=( (not A236)  and  (not A235) );
 a40335a <=( (not A268)  and  (not A267) );
 a40336a <=( a40335a  and  a40332a );
 a40339a <=( (not A298)  and  (not A269) );
 a40342a <=( (not A301)  and  (not A299) );
 a40343a <=( a40342a  and  a40339a );
 a40344a <=( a40343a  and  a40336a );
 a40348a <=( A166  and  (not A167) );
 a40349a <=( A170  and  a40348a );
 a40352a <=( (not A200)  and  (not A199) );
 a40355a <=( (not A234)  and  (not A202) );
 a40356a <=( a40355a  and  a40352a );
 a40357a <=( a40356a  and  a40349a );
 a40360a <=( (not A236)  and  (not A235) );
 a40363a <=( (not A266)  and  (not A265) );
 a40364a <=( a40363a  and  a40360a );
 a40367a <=( (not A300)  and  (not A268) );
 a40370a <=( (not A302)  and  (not A301) );
 a40371a <=( a40370a  and  a40367a );
 a40372a <=( a40371a  and  a40364a );
 a40376a <=( A166  and  (not A167) );
 a40377a <=( A170  and  a40376a );
 a40380a <=( (not A200)  and  (not A199) );
 a40383a <=( (not A234)  and  (not A202) );
 a40384a <=( a40383a  and  a40380a );
 a40385a <=( a40384a  and  a40377a );
 a40388a <=( (not A236)  and  (not A235) );
 a40391a <=( (not A266)  and  (not A265) );
 a40392a <=( a40391a  and  a40388a );
 a40395a <=( (not A298)  and  (not A268) );
 a40398a <=( (not A301)  and  (not A299) );
 a40399a <=( a40398a  and  a40395a );
 a40400a <=( a40399a  and  a40392a );
 a40404a <=( A166  and  (not A167) );
 a40405a <=( A170  and  a40404a );
 a40408a <=( (not A200)  and  (not A199) );
 a40411a <=( (not A232)  and  (not A202) );
 a40412a <=( a40411a  and  a40408a );
 a40413a <=( a40412a  and  a40405a );
 a40416a <=( (not A235)  and  (not A233) );
 a40419a <=( (not A268)  and  (not A267) );
 a40420a <=( a40419a  and  a40416a );
 a40423a <=( (not A300)  and  (not A269) );
 a40426a <=( (not A302)  and  (not A301) );
 a40427a <=( a40426a  and  a40423a );
 a40428a <=( a40427a  and  a40420a );
 a40432a <=( A166  and  (not A167) );
 a40433a <=( A170  and  a40432a );
 a40436a <=( (not A200)  and  (not A199) );
 a40439a <=( (not A232)  and  (not A202) );
 a40440a <=( a40439a  and  a40436a );
 a40441a <=( a40440a  and  a40433a );
 a40444a <=( (not A235)  and  (not A233) );
 a40447a <=( (not A268)  and  (not A267) );
 a40448a <=( a40447a  and  a40444a );
 a40451a <=( (not A298)  and  (not A269) );
 a40454a <=( (not A301)  and  (not A299) );
 a40455a <=( a40454a  and  a40451a );
 a40456a <=( a40455a  and  a40448a );
 a40460a <=( A166  and  (not A167) );
 a40461a <=( A170  and  a40460a );
 a40464a <=( (not A200)  and  (not A199) );
 a40467a <=( (not A232)  and  (not A202) );
 a40468a <=( a40467a  and  a40464a );
 a40469a <=( a40468a  and  a40461a );
 a40472a <=( (not A235)  and  (not A233) );
 a40475a <=( (not A266)  and  (not A265) );
 a40476a <=( a40475a  and  a40472a );
 a40479a <=( (not A300)  and  (not A268) );
 a40482a <=( (not A302)  and  (not A301) );
 a40483a <=( a40482a  and  a40479a );
 a40484a <=( a40483a  and  a40476a );
 a40488a <=( A166  and  (not A167) );
 a40489a <=( A170  and  a40488a );
 a40492a <=( (not A200)  and  (not A199) );
 a40495a <=( (not A232)  and  (not A202) );
 a40496a <=( a40495a  and  a40492a );
 a40497a <=( a40496a  and  a40489a );
 a40500a <=( (not A235)  and  (not A233) );
 a40503a <=( (not A266)  and  (not A265) );
 a40504a <=( a40503a  and  a40500a );
 a40507a <=( (not A298)  and  (not A268) );
 a40510a <=( (not A301)  and  (not A299) );
 a40511a <=( a40510a  and  a40507a );
 a40512a <=( a40511a  and  a40504a );
 a40516a <=( (not A202)  and  (not A201) );
 a40517a <=( A169  and  a40516a );
 a40520a <=( (not A234)  and  (not A203) );
 a40523a <=( (not A236)  and  (not A235) );
 a40524a <=( a40523a  and  a40520a );
 a40525a <=( a40524a  and  a40517a );
 a40528a <=( A266  and  A265 );
 a40531a <=( (not A268)  and  (not A267) );
 a40532a <=( a40531a  and  a40528a );
 a40535a <=( A299  and  A298 );
 a40538a <=( (not A301)  and  (not A300) );
 a40539a <=( a40538a  and  a40535a );
 a40540a <=( a40539a  and  a40532a );
 a40544a <=( (not A202)  and  (not A201) );
 a40545a <=( A169  and  a40544a );
 a40548a <=( A232  and  (not A203) );
 a40551a <=( (not A234)  and  A233 );
 a40552a <=( a40551a  and  a40548a );
 a40553a <=( a40552a  and  a40545a );
 a40556a <=( (not A267)  and  (not A235) );
 a40559a <=( (not A269)  and  (not A268) );
 a40560a <=( a40559a  and  a40556a );
 a40563a <=( A299  and  A298 );
 a40566a <=( (not A301)  and  (not A300) );
 a40567a <=( a40566a  and  a40563a );
 a40568a <=( a40567a  and  a40560a );
 a40572a <=( (not A202)  and  (not A201) );
 a40573a <=( A169  and  a40572a );
 a40576a <=( A232  and  (not A203) );
 a40579a <=( (not A234)  and  A233 );
 a40580a <=( a40579a  and  a40576a );
 a40581a <=( a40580a  and  a40573a );
 a40584a <=( A265  and  (not A235) );
 a40587a <=( (not A267)  and  A266 );
 a40588a <=( a40587a  and  a40584a );
 a40591a <=( (not A300)  and  (not A268) );
 a40594a <=( (not A302)  and  (not A301) );
 a40595a <=( a40594a  and  a40591a );
 a40596a <=( a40595a  and  a40588a );
 a40600a <=( (not A202)  and  (not A201) );
 a40601a <=( A169  and  a40600a );
 a40604a <=( A232  and  (not A203) );
 a40607a <=( (not A234)  and  A233 );
 a40608a <=( a40607a  and  a40604a );
 a40609a <=( a40608a  and  a40601a );
 a40612a <=( A265  and  (not A235) );
 a40615a <=( (not A267)  and  A266 );
 a40616a <=( a40615a  and  a40612a );
 a40619a <=( (not A298)  and  (not A268) );
 a40622a <=( (not A301)  and  (not A299) );
 a40623a <=( a40622a  and  a40619a );
 a40624a <=( a40623a  and  a40616a );
 a40628a <=( (not A202)  and  (not A201) );
 a40629a <=( A169  and  a40628a );
 a40632a <=( A232  and  (not A203) );
 a40635a <=( (not A234)  and  A233 );
 a40636a <=( a40635a  and  a40632a );
 a40637a <=( a40636a  and  a40629a );
 a40640a <=( (not A265)  and  (not A235) );
 a40643a <=( (not A268)  and  (not A266) );
 a40644a <=( a40643a  and  a40640a );
 a40647a <=( A299  and  A298 );
 a40650a <=( (not A301)  and  (not A300) );
 a40651a <=( a40650a  and  a40647a );
 a40652a <=( a40651a  and  a40644a );
 a40656a <=( (not A202)  and  (not A201) );
 a40657a <=( A169  and  a40656a );
 a40660a <=( (not A232)  and  (not A203) );
 a40663a <=( (not A235)  and  (not A233) );
 a40664a <=( a40663a  and  a40660a );
 a40665a <=( a40664a  and  a40657a );
 a40668a <=( A266  and  A265 );
 a40671a <=( (not A268)  and  (not A267) );
 a40672a <=( a40671a  and  a40668a );
 a40675a <=( A299  and  A298 );
 a40678a <=( (not A301)  and  (not A300) );
 a40679a <=( a40678a  and  a40675a );
 a40680a <=( a40679a  and  a40672a );
 a40684a <=( A200  and  A199 );
 a40685a <=( A169  and  a40684a );
 a40688a <=( (not A202)  and  (not A201) );
 a40691a <=( (not A235)  and  (not A234) );
 a40692a <=( a40691a  and  a40688a );
 a40693a <=( a40692a  and  a40685a );
 a40696a <=( (not A267)  and  (not A236) );
 a40699a <=( (not A269)  and  (not A268) );
 a40700a <=( a40699a  and  a40696a );
 a40703a <=( A299  and  A298 );
 a40706a <=( (not A301)  and  (not A300) );
 a40707a <=( a40706a  and  a40703a );
 a40708a <=( a40707a  and  a40700a );
 a40712a <=( A200  and  A199 );
 a40713a <=( A169  and  a40712a );
 a40716a <=( (not A202)  and  (not A201) );
 a40719a <=( (not A235)  and  (not A234) );
 a40720a <=( a40719a  and  a40716a );
 a40721a <=( a40720a  and  a40713a );
 a40724a <=( A265  and  (not A236) );
 a40727a <=( (not A267)  and  A266 );
 a40728a <=( a40727a  and  a40724a );
 a40731a <=( (not A300)  and  (not A268) );
 a40734a <=( (not A302)  and  (not A301) );
 a40735a <=( a40734a  and  a40731a );
 a40736a <=( a40735a  and  a40728a );
 a40740a <=( A200  and  A199 );
 a40741a <=( A169  and  a40740a );
 a40744a <=( (not A202)  and  (not A201) );
 a40747a <=( (not A235)  and  (not A234) );
 a40748a <=( a40747a  and  a40744a );
 a40749a <=( a40748a  and  a40741a );
 a40752a <=( A265  and  (not A236) );
 a40755a <=( (not A267)  and  A266 );
 a40756a <=( a40755a  and  a40752a );
 a40759a <=( (not A298)  and  (not A268) );
 a40762a <=( (not A301)  and  (not A299) );
 a40763a <=( a40762a  and  a40759a );
 a40764a <=( a40763a  and  a40756a );
 a40768a <=( A200  and  A199 );
 a40769a <=( A169  and  a40768a );
 a40772a <=( (not A202)  and  (not A201) );
 a40775a <=( (not A235)  and  (not A234) );
 a40776a <=( a40775a  and  a40772a );
 a40777a <=( a40776a  and  a40769a );
 a40780a <=( (not A265)  and  (not A236) );
 a40783a <=( (not A268)  and  (not A266) );
 a40784a <=( a40783a  and  a40780a );
 a40787a <=( A299  and  A298 );
 a40790a <=( (not A301)  and  (not A300) );
 a40791a <=( a40790a  and  a40787a );
 a40792a <=( a40791a  and  a40784a );
 a40796a <=( A200  and  A199 );
 a40797a <=( A169  and  a40796a );
 a40800a <=( (not A202)  and  (not A201) );
 a40803a <=( A233  and  A232 );
 a40804a <=( a40803a  and  a40800a );
 a40805a <=( a40804a  and  a40797a );
 a40808a <=( (not A235)  and  (not A234) );
 a40811a <=( (not A268)  and  (not A267) );
 a40812a <=( a40811a  and  a40808a );
 a40815a <=( (not A300)  and  (not A269) );
 a40818a <=( (not A302)  and  (not A301) );
 a40819a <=( a40818a  and  a40815a );
 a40820a <=( a40819a  and  a40812a );
 a40824a <=( A200  and  A199 );
 a40825a <=( A169  and  a40824a );
 a40828a <=( (not A202)  and  (not A201) );
 a40831a <=( A233  and  A232 );
 a40832a <=( a40831a  and  a40828a );
 a40833a <=( a40832a  and  a40825a );
 a40836a <=( (not A235)  and  (not A234) );
 a40839a <=( (not A268)  and  (not A267) );
 a40840a <=( a40839a  and  a40836a );
 a40843a <=( (not A298)  and  (not A269) );
 a40846a <=( (not A301)  and  (not A299) );
 a40847a <=( a40846a  and  a40843a );
 a40848a <=( a40847a  and  a40840a );
 a40852a <=( A200  and  A199 );
 a40853a <=( A169  and  a40852a );
 a40856a <=( (not A202)  and  (not A201) );
 a40859a <=( A233  and  A232 );
 a40860a <=( a40859a  and  a40856a );
 a40861a <=( a40860a  and  a40853a );
 a40864a <=( (not A235)  and  (not A234) );
 a40867a <=( (not A266)  and  (not A265) );
 a40868a <=( a40867a  and  a40864a );
 a40871a <=( (not A300)  and  (not A268) );
 a40874a <=( (not A302)  and  (not A301) );
 a40875a <=( a40874a  and  a40871a );
 a40876a <=( a40875a  and  a40868a );
 a40880a <=( A200  and  A199 );
 a40881a <=( A169  and  a40880a );
 a40884a <=( (not A202)  and  (not A201) );
 a40887a <=( A233  and  A232 );
 a40888a <=( a40887a  and  a40884a );
 a40889a <=( a40888a  and  a40881a );
 a40892a <=( (not A235)  and  (not A234) );
 a40895a <=( (not A266)  and  (not A265) );
 a40896a <=( a40895a  and  a40892a );
 a40899a <=( (not A298)  and  (not A268) );
 a40902a <=( (not A301)  and  (not A299) );
 a40903a <=( a40902a  and  a40899a );
 a40904a <=( a40903a  and  a40896a );
 a40908a <=( A200  and  A199 );
 a40909a <=( A169  and  a40908a );
 a40912a <=( (not A202)  and  (not A201) );
 a40915a <=( (not A233)  and  (not A232) );
 a40916a <=( a40915a  and  a40912a );
 a40917a <=( a40916a  and  a40909a );
 a40920a <=( (not A267)  and  (not A235) );
 a40923a <=( (not A269)  and  (not A268) );
 a40924a <=( a40923a  and  a40920a );
 a40927a <=( A299  and  A298 );
 a40930a <=( (not A301)  and  (not A300) );
 a40931a <=( a40930a  and  a40927a );
 a40932a <=( a40931a  and  a40924a );
 a40936a <=( A200  and  A199 );
 a40937a <=( A169  and  a40936a );
 a40940a <=( (not A202)  and  (not A201) );
 a40943a <=( (not A233)  and  (not A232) );
 a40944a <=( a40943a  and  a40940a );
 a40945a <=( a40944a  and  a40937a );
 a40948a <=( A265  and  (not A235) );
 a40951a <=( (not A267)  and  A266 );
 a40952a <=( a40951a  and  a40948a );
 a40955a <=( (not A300)  and  (not A268) );
 a40958a <=( (not A302)  and  (not A301) );
 a40959a <=( a40958a  and  a40955a );
 a40960a <=( a40959a  and  a40952a );
 a40964a <=( A200  and  A199 );
 a40965a <=( A169  and  a40964a );
 a40968a <=( (not A202)  and  (not A201) );
 a40971a <=( (not A233)  and  (not A232) );
 a40972a <=( a40971a  and  a40968a );
 a40973a <=( a40972a  and  a40965a );
 a40976a <=( A265  and  (not A235) );
 a40979a <=( (not A267)  and  A266 );
 a40980a <=( a40979a  and  a40976a );
 a40983a <=( (not A298)  and  (not A268) );
 a40986a <=( (not A301)  and  (not A299) );
 a40987a <=( a40986a  and  a40983a );
 a40988a <=( a40987a  and  a40980a );
 a40992a <=( A200  and  A199 );
 a40993a <=( A169  and  a40992a );
 a40996a <=( (not A202)  and  (not A201) );
 a40999a <=( (not A233)  and  (not A232) );
 a41000a <=( a40999a  and  a40996a );
 a41001a <=( a41000a  and  a40993a );
 a41004a <=( (not A265)  and  (not A235) );
 a41007a <=( (not A268)  and  (not A266) );
 a41008a <=( a41007a  and  a41004a );
 a41011a <=( A299  and  A298 );
 a41014a <=( (not A301)  and  (not A300) );
 a41015a <=( a41014a  and  a41011a );
 a41016a <=( a41015a  and  a41008a );
 a41020a <=( (not A200)  and  (not A199) );
 a41021a <=( A169  and  a41020a );
 a41024a <=( (not A234)  and  (not A202) );
 a41027a <=( (not A236)  and  (not A235) );
 a41028a <=( a41027a  and  a41024a );
 a41029a <=( a41028a  and  a41021a );
 a41032a <=( A266  and  A265 );
 a41035a <=( (not A268)  and  (not A267) );
 a41036a <=( a41035a  and  a41032a );
 a41039a <=( A299  and  A298 );
 a41042a <=( (not A301)  and  (not A300) );
 a41043a <=( a41042a  and  a41039a );
 a41044a <=( a41043a  and  a41036a );
 a41048a <=( (not A200)  and  (not A199) );
 a41049a <=( A169  and  a41048a );
 a41052a <=( A232  and  (not A202) );
 a41055a <=( (not A234)  and  A233 );
 a41056a <=( a41055a  and  a41052a );
 a41057a <=( a41056a  and  a41049a );
 a41060a <=( (not A267)  and  (not A235) );
 a41063a <=( (not A269)  and  (not A268) );
 a41064a <=( a41063a  and  a41060a );
 a41067a <=( A299  and  A298 );
 a41070a <=( (not A301)  and  (not A300) );
 a41071a <=( a41070a  and  a41067a );
 a41072a <=( a41071a  and  a41064a );
 a41076a <=( (not A200)  and  (not A199) );
 a41077a <=( A169  and  a41076a );
 a41080a <=( A232  and  (not A202) );
 a41083a <=( (not A234)  and  A233 );
 a41084a <=( a41083a  and  a41080a );
 a41085a <=( a41084a  and  a41077a );
 a41088a <=( A265  and  (not A235) );
 a41091a <=( (not A267)  and  A266 );
 a41092a <=( a41091a  and  a41088a );
 a41095a <=( (not A300)  and  (not A268) );
 a41098a <=( (not A302)  and  (not A301) );
 a41099a <=( a41098a  and  a41095a );
 a41100a <=( a41099a  and  a41092a );
 a41104a <=( (not A200)  and  (not A199) );
 a41105a <=( A169  and  a41104a );
 a41108a <=( A232  and  (not A202) );
 a41111a <=( (not A234)  and  A233 );
 a41112a <=( a41111a  and  a41108a );
 a41113a <=( a41112a  and  a41105a );
 a41116a <=( A265  and  (not A235) );
 a41119a <=( (not A267)  and  A266 );
 a41120a <=( a41119a  and  a41116a );
 a41123a <=( (not A298)  and  (not A268) );
 a41126a <=( (not A301)  and  (not A299) );
 a41127a <=( a41126a  and  a41123a );
 a41128a <=( a41127a  and  a41120a );
 a41132a <=( (not A200)  and  (not A199) );
 a41133a <=( A169  and  a41132a );
 a41136a <=( A232  and  (not A202) );
 a41139a <=( (not A234)  and  A233 );
 a41140a <=( a41139a  and  a41136a );
 a41141a <=( a41140a  and  a41133a );
 a41144a <=( (not A265)  and  (not A235) );
 a41147a <=( (not A268)  and  (not A266) );
 a41148a <=( a41147a  and  a41144a );
 a41151a <=( A299  and  A298 );
 a41154a <=( (not A301)  and  (not A300) );
 a41155a <=( a41154a  and  a41151a );
 a41156a <=( a41155a  and  a41148a );
 a41160a <=( (not A200)  and  (not A199) );
 a41161a <=( A169  and  a41160a );
 a41164a <=( (not A232)  and  (not A202) );
 a41167a <=( (not A235)  and  (not A233) );
 a41168a <=( a41167a  and  a41164a );
 a41169a <=( a41168a  and  a41161a );
 a41172a <=( A266  and  A265 );
 a41175a <=( (not A268)  and  (not A267) );
 a41176a <=( a41175a  and  a41172a );
 a41179a <=( A299  and  A298 );
 a41182a <=( (not A301)  and  (not A300) );
 a41183a <=( a41182a  and  a41179a );
 a41184a <=( a41183a  and  a41176a );
 a41188a <=( (not A166)  and  (not A167) );
 a41189a <=( (not A169)  and  a41188a );
 a41192a <=( (not A234)  and  A202 );
 a41195a <=( (not A236)  and  (not A235) );
 a41196a <=( a41195a  and  a41192a );
 a41197a <=( a41196a  and  a41189a );
 a41200a <=( A266  and  A265 );
 a41203a <=( (not A268)  and  (not A267) );
 a41204a <=( a41203a  and  a41200a );
 a41207a <=( A299  and  A298 );
 a41210a <=( (not A301)  and  (not A300) );
 a41211a <=( a41210a  and  a41207a );
 a41212a <=( a41211a  and  a41204a );
 a41216a <=( (not A166)  and  (not A167) );
 a41217a <=( (not A169)  and  a41216a );
 a41220a <=( A232  and  A202 );
 a41223a <=( (not A234)  and  A233 );
 a41224a <=( a41223a  and  a41220a );
 a41225a <=( a41224a  and  a41217a );
 a41228a <=( (not A267)  and  (not A235) );
 a41231a <=( (not A269)  and  (not A268) );
 a41232a <=( a41231a  and  a41228a );
 a41235a <=( A299  and  A298 );
 a41238a <=( (not A301)  and  (not A300) );
 a41239a <=( a41238a  and  a41235a );
 a41240a <=( a41239a  and  a41232a );
 a41244a <=( (not A166)  and  (not A167) );
 a41245a <=( (not A169)  and  a41244a );
 a41248a <=( A232  and  A202 );
 a41251a <=( (not A234)  and  A233 );
 a41252a <=( a41251a  and  a41248a );
 a41253a <=( a41252a  and  a41245a );
 a41256a <=( A265  and  (not A235) );
 a41259a <=( (not A267)  and  A266 );
 a41260a <=( a41259a  and  a41256a );
 a41263a <=( (not A300)  and  (not A268) );
 a41266a <=( (not A302)  and  (not A301) );
 a41267a <=( a41266a  and  a41263a );
 a41268a <=( a41267a  and  a41260a );
 a41272a <=( (not A166)  and  (not A167) );
 a41273a <=( (not A169)  and  a41272a );
 a41276a <=( A232  and  A202 );
 a41279a <=( (not A234)  and  A233 );
 a41280a <=( a41279a  and  a41276a );
 a41281a <=( a41280a  and  a41273a );
 a41284a <=( A265  and  (not A235) );
 a41287a <=( (not A267)  and  A266 );
 a41288a <=( a41287a  and  a41284a );
 a41291a <=( (not A298)  and  (not A268) );
 a41294a <=( (not A301)  and  (not A299) );
 a41295a <=( a41294a  and  a41291a );
 a41296a <=( a41295a  and  a41288a );
 a41300a <=( (not A166)  and  (not A167) );
 a41301a <=( (not A169)  and  a41300a );
 a41304a <=( A232  and  A202 );
 a41307a <=( (not A234)  and  A233 );
 a41308a <=( a41307a  and  a41304a );
 a41309a <=( a41308a  and  a41301a );
 a41312a <=( (not A265)  and  (not A235) );
 a41315a <=( (not A268)  and  (not A266) );
 a41316a <=( a41315a  and  a41312a );
 a41319a <=( A299  and  A298 );
 a41322a <=( (not A301)  and  (not A300) );
 a41323a <=( a41322a  and  a41319a );
 a41324a <=( a41323a  and  a41316a );
 a41328a <=( (not A166)  and  (not A167) );
 a41329a <=( (not A169)  and  a41328a );
 a41332a <=( (not A232)  and  A202 );
 a41335a <=( (not A235)  and  (not A233) );
 a41336a <=( a41335a  and  a41332a );
 a41337a <=( a41336a  and  a41329a );
 a41340a <=( A266  and  A265 );
 a41343a <=( (not A268)  and  (not A267) );
 a41344a <=( a41343a  and  a41340a );
 a41347a <=( A299  and  A298 );
 a41350a <=( (not A301)  and  (not A300) );
 a41351a <=( a41350a  and  a41347a );
 a41352a <=( a41351a  and  a41344a );
 a41356a <=( (not A166)  and  (not A167) );
 a41357a <=( (not A169)  and  a41356a );
 a41360a <=( A201  and  A199 );
 a41363a <=( (not A235)  and  (not A234) );
 a41364a <=( a41363a  and  a41360a );
 a41365a <=( a41364a  and  a41357a );
 a41368a <=( (not A267)  and  (not A236) );
 a41371a <=( (not A269)  and  (not A268) );
 a41372a <=( a41371a  and  a41368a );
 a41375a <=( A299  and  A298 );
 a41378a <=( (not A301)  and  (not A300) );
 a41379a <=( a41378a  and  a41375a );
 a41380a <=( a41379a  and  a41372a );
 a41384a <=( (not A166)  and  (not A167) );
 a41385a <=( (not A169)  and  a41384a );
 a41388a <=( A201  and  A199 );
 a41391a <=( (not A235)  and  (not A234) );
 a41392a <=( a41391a  and  a41388a );
 a41393a <=( a41392a  and  a41385a );
 a41396a <=( A265  and  (not A236) );
 a41399a <=( (not A267)  and  A266 );
 a41400a <=( a41399a  and  a41396a );
 a41403a <=( (not A300)  and  (not A268) );
 a41406a <=( (not A302)  and  (not A301) );
 a41407a <=( a41406a  and  a41403a );
 a41408a <=( a41407a  and  a41400a );
 a41412a <=( (not A166)  and  (not A167) );
 a41413a <=( (not A169)  and  a41412a );
 a41416a <=( A201  and  A199 );
 a41419a <=( (not A235)  and  (not A234) );
 a41420a <=( a41419a  and  a41416a );
 a41421a <=( a41420a  and  a41413a );
 a41424a <=( A265  and  (not A236) );
 a41427a <=( (not A267)  and  A266 );
 a41428a <=( a41427a  and  a41424a );
 a41431a <=( (not A298)  and  (not A268) );
 a41434a <=( (not A301)  and  (not A299) );
 a41435a <=( a41434a  and  a41431a );
 a41436a <=( a41435a  and  a41428a );
 a41440a <=( (not A166)  and  (not A167) );
 a41441a <=( (not A169)  and  a41440a );
 a41444a <=( A201  and  A199 );
 a41447a <=( (not A235)  and  (not A234) );
 a41448a <=( a41447a  and  a41444a );
 a41449a <=( a41448a  and  a41441a );
 a41452a <=( (not A265)  and  (not A236) );
 a41455a <=( (not A268)  and  (not A266) );
 a41456a <=( a41455a  and  a41452a );
 a41459a <=( A299  and  A298 );
 a41462a <=( (not A301)  and  (not A300) );
 a41463a <=( a41462a  and  a41459a );
 a41464a <=( a41463a  and  a41456a );
 a41468a <=( (not A166)  and  (not A167) );
 a41469a <=( (not A169)  and  a41468a );
 a41472a <=( A201  and  A199 );
 a41475a <=( A233  and  A232 );
 a41476a <=( a41475a  and  a41472a );
 a41477a <=( a41476a  and  a41469a );
 a41480a <=( (not A235)  and  (not A234) );
 a41483a <=( (not A268)  and  (not A267) );
 a41484a <=( a41483a  and  a41480a );
 a41487a <=( (not A300)  and  (not A269) );
 a41490a <=( (not A302)  and  (not A301) );
 a41491a <=( a41490a  and  a41487a );
 a41492a <=( a41491a  and  a41484a );
 a41496a <=( (not A166)  and  (not A167) );
 a41497a <=( (not A169)  and  a41496a );
 a41500a <=( A201  and  A199 );
 a41503a <=( A233  and  A232 );
 a41504a <=( a41503a  and  a41500a );
 a41505a <=( a41504a  and  a41497a );
 a41508a <=( (not A235)  and  (not A234) );
 a41511a <=( (not A268)  and  (not A267) );
 a41512a <=( a41511a  and  a41508a );
 a41515a <=( (not A298)  and  (not A269) );
 a41518a <=( (not A301)  and  (not A299) );
 a41519a <=( a41518a  and  a41515a );
 a41520a <=( a41519a  and  a41512a );
 a41524a <=( (not A166)  and  (not A167) );
 a41525a <=( (not A169)  and  a41524a );
 a41528a <=( A201  and  A199 );
 a41531a <=( A233  and  A232 );
 a41532a <=( a41531a  and  a41528a );
 a41533a <=( a41532a  and  a41525a );
 a41536a <=( (not A235)  and  (not A234) );
 a41539a <=( (not A266)  and  (not A265) );
 a41540a <=( a41539a  and  a41536a );
 a41543a <=( (not A300)  and  (not A268) );
 a41546a <=( (not A302)  and  (not A301) );
 a41547a <=( a41546a  and  a41543a );
 a41548a <=( a41547a  and  a41540a );
 a41552a <=( (not A166)  and  (not A167) );
 a41553a <=( (not A169)  and  a41552a );
 a41556a <=( A201  and  A199 );
 a41559a <=( A233  and  A232 );
 a41560a <=( a41559a  and  a41556a );
 a41561a <=( a41560a  and  a41553a );
 a41564a <=( (not A235)  and  (not A234) );
 a41567a <=( (not A266)  and  (not A265) );
 a41568a <=( a41567a  and  a41564a );
 a41571a <=( (not A298)  and  (not A268) );
 a41574a <=( (not A301)  and  (not A299) );
 a41575a <=( a41574a  and  a41571a );
 a41576a <=( a41575a  and  a41568a );
 a41580a <=( (not A166)  and  (not A167) );
 a41581a <=( (not A169)  and  a41580a );
 a41584a <=( A201  and  A199 );
 a41587a <=( (not A233)  and  (not A232) );
 a41588a <=( a41587a  and  a41584a );
 a41589a <=( a41588a  and  a41581a );
 a41592a <=( (not A267)  and  (not A235) );
 a41595a <=( (not A269)  and  (not A268) );
 a41596a <=( a41595a  and  a41592a );
 a41599a <=( A299  and  A298 );
 a41602a <=( (not A301)  and  (not A300) );
 a41603a <=( a41602a  and  a41599a );
 a41604a <=( a41603a  and  a41596a );
 a41608a <=( (not A166)  and  (not A167) );
 a41609a <=( (not A169)  and  a41608a );
 a41612a <=( A201  and  A199 );
 a41615a <=( (not A233)  and  (not A232) );
 a41616a <=( a41615a  and  a41612a );
 a41617a <=( a41616a  and  a41609a );
 a41620a <=( A265  and  (not A235) );
 a41623a <=( (not A267)  and  A266 );
 a41624a <=( a41623a  and  a41620a );
 a41627a <=( (not A300)  and  (not A268) );
 a41630a <=( (not A302)  and  (not A301) );
 a41631a <=( a41630a  and  a41627a );
 a41632a <=( a41631a  and  a41624a );
 a41636a <=( (not A166)  and  (not A167) );
 a41637a <=( (not A169)  and  a41636a );
 a41640a <=( A201  and  A199 );
 a41643a <=( (not A233)  and  (not A232) );
 a41644a <=( a41643a  and  a41640a );
 a41645a <=( a41644a  and  a41637a );
 a41648a <=( A265  and  (not A235) );
 a41651a <=( (not A267)  and  A266 );
 a41652a <=( a41651a  and  a41648a );
 a41655a <=( (not A298)  and  (not A268) );
 a41658a <=( (not A301)  and  (not A299) );
 a41659a <=( a41658a  and  a41655a );
 a41660a <=( a41659a  and  a41652a );
 a41664a <=( (not A166)  and  (not A167) );
 a41665a <=( (not A169)  and  a41664a );
 a41668a <=( A201  and  A199 );
 a41671a <=( (not A233)  and  (not A232) );
 a41672a <=( a41671a  and  a41668a );
 a41673a <=( a41672a  and  a41665a );
 a41676a <=( (not A265)  and  (not A235) );
 a41679a <=( (not A268)  and  (not A266) );
 a41680a <=( a41679a  and  a41676a );
 a41683a <=( A299  and  A298 );
 a41686a <=( (not A301)  and  (not A300) );
 a41687a <=( a41686a  and  a41683a );
 a41688a <=( a41687a  and  a41680a );
 a41692a <=( (not A166)  and  (not A167) );
 a41693a <=( (not A169)  and  a41692a );
 a41696a <=( A201  and  A200 );
 a41699a <=( (not A235)  and  (not A234) );
 a41700a <=( a41699a  and  a41696a );
 a41701a <=( a41700a  and  a41693a );
 a41704a <=( (not A267)  and  (not A236) );
 a41707a <=( (not A269)  and  (not A268) );
 a41708a <=( a41707a  and  a41704a );
 a41711a <=( A299  and  A298 );
 a41714a <=( (not A301)  and  (not A300) );
 a41715a <=( a41714a  and  a41711a );
 a41716a <=( a41715a  and  a41708a );
 a41720a <=( (not A166)  and  (not A167) );
 a41721a <=( (not A169)  and  a41720a );
 a41724a <=( A201  and  A200 );
 a41727a <=( (not A235)  and  (not A234) );
 a41728a <=( a41727a  and  a41724a );
 a41729a <=( a41728a  and  a41721a );
 a41732a <=( A265  and  (not A236) );
 a41735a <=( (not A267)  and  A266 );
 a41736a <=( a41735a  and  a41732a );
 a41739a <=( (not A300)  and  (not A268) );
 a41742a <=( (not A302)  and  (not A301) );
 a41743a <=( a41742a  and  a41739a );
 a41744a <=( a41743a  and  a41736a );
 a41748a <=( (not A166)  and  (not A167) );
 a41749a <=( (not A169)  and  a41748a );
 a41752a <=( A201  and  A200 );
 a41755a <=( (not A235)  and  (not A234) );
 a41756a <=( a41755a  and  a41752a );
 a41757a <=( a41756a  and  a41749a );
 a41760a <=( A265  and  (not A236) );
 a41763a <=( (not A267)  and  A266 );
 a41764a <=( a41763a  and  a41760a );
 a41767a <=( (not A298)  and  (not A268) );
 a41770a <=( (not A301)  and  (not A299) );
 a41771a <=( a41770a  and  a41767a );
 a41772a <=( a41771a  and  a41764a );
 a41776a <=( (not A166)  and  (not A167) );
 a41777a <=( (not A169)  and  a41776a );
 a41780a <=( A201  and  A200 );
 a41783a <=( (not A235)  and  (not A234) );
 a41784a <=( a41783a  and  a41780a );
 a41785a <=( a41784a  and  a41777a );
 a41788a <=( (not A265)  and  (not A236) );
 a41791a <=( (not A268)  and  (not A266) );
 a41792a <=( a41791a  and  a41788a );
 a41795a <=( A299  and  A298 );
 a41798a <=( (not A301)  and  (not A300) );
 a41799a <=( a41798a  and  a41795a );
 a41800a <=( a41799a  and  a41792a );
 a41804a <=( (not A166)  and  (not A167) );
 a41805a <=( (not A169)  and  a41804a );
 a41808a <=( A201  and  A200 );
 a41811a <=( A233  and  A232 );
 a41812a <=( a41811a  and  a41808a );
 a41813a <=( a41812a  and  a41805a );
 a41816a <=( (not A235)  and  (not A234) );
 a41819a <=( (not A268)  and  (not A267) );
 a41820a <=( a41819a  and  a41816a );
 a41823a <=( (not A300)  and  (not A269) );
 a41826a <=( (not A302)  and  (not A301) );
 a41827a <=( a41826a  and  a41823a );
 a41828a <=( a41827a  and  a41820a );
 a41832a <=( (not A166)  and  (not A167) );
 a41833a <=( (not A169)  and  a41832a );
 a41836a <=( A201  and  A200 );
 a41839a <=( A233  and  A232 );
 a41840a <=( a41839a  and  a41836a );
 a41841a <=( a41840a  and  a41833a );
 a41844a <=( (not A235)  and  (not A234) );
 a41847a <=( (not A268)  and  (not A267) );
 a41848a <=( a41847a  and  a41844a );
 a41851a <=( (not A298)  and  (not A269) );
 a41854a <=( (not A301)  and  (not A299) );
 a41855a <=( a41854a  and  a41851a );
 a41856a <=( a41855a  and  a41848a );
 a41860a <=( (not A166)  and  (not A167) );
 a41861a <=( (not A169)  and  a41860a );
 a41864a <=( A201  and  A200 );
 a41867a <=( A233  and  A232 );
 a41868a <=( a41867a  and  a41864a );
 a41869a <=( a41868a  and  a41861a );
 a41872a <=( (not A235)  and  (not A234) );
 a41875a <=( (not A266)  and  (not A265) );
 a41876a <=( a41875a  and  a41872a );
 a41879a <=( (not A300)  and  (not A268) );
 a41882a <=( (not A302)  and  (not A301) );
 a41883a <=( a41882a  and  a41879a );
 a41884a <=( a41883a  and  a41876a );
 a41888a <=( (not A166)  and  (not A167) );
 a41889a <=( (not A169)  and  a41888a );
 a41892a <=( A201  and  A200 );
 a41895a <=( A233  and  A232 );
 a41896a <=( a41895a  and  a41892a );
 a41897a <=( a41896a  and  a41889a );
 a41900a <=( (not A235)  and  (not A234) );
 a41903a <=( (not A266)  and  (not A265) );
 a41904a <=( a41903a  and  a41900a );
 a41907a <=( (not A298)  and  (not A268) );
 a41910a <=( (not A301)  and  (not A299) );
 a41911a <=( a41910a  and  a41907a );
 a41912a <=( a41911a  and  a41904a );
 a41916a <=( (not A166)  and  (not A167) );
 a41917a <=( (not A169)  and  a41916a );
 a41920a <=( A201  and  A200 );
 a41923a <=( (not A233)  and  (not A232) );
 a41924a <=( a41923a  and  a41920a );
 a41925a <=( a41924a  and  a41917a );
 a41928a <=( (not A267)  and  (not A235) );
 a41931a <=( (not A269)  and  (not A268) );
 a41932a <=( a41931a  and  a41928a );
 a41935a <=( A299  and  A298 );
 a41938a <=( (not A301)  and  (not A300) );
 a41939a <=( a41938a  and  a41935a );
 a41940a <=( a41939a  and  a41932a );
 a41944a <=( (not A166)  and  (not A167) );
 a41945a <=( (not A169)  and  a41944a );
 a41948a <=( A201  and  A200 );
 a41951a <=( (not A233)  and  (not A232) );
 a41952a <=( a41951a  and  a41948a );
 a41953a <=( a41952a  and  a41945a );
 a41956a <=( A265  and  (not A235) );
 a41959a <=( (not A267)  and  A266 );
 a41960a <=( a41959a  and  a41956a );
 a41963a <=( (not A300)  and  (not A268) );
 a41966a <=( (not A302)  and  (not A301) );
 a41967a <=( a41966a  and  a41963a );
 a41968a <=( a41967a  and  a41960a );
 a41972a <=( (not A166)  and  (not A167) );
 a41973a <=( (not A169)  and  a41972a );
 a41976a <=( A201  and  A200 );
 a41979a <=( (not A233)  and  (not A232) );
 a41980a <=( a41979a  and  a41976a );
 a41981a <=( a41980a  and  a41973a );
 a41984a <=( A265  and  (not A235) );
 a41987a <=( (not A267)  and  A266 );
 a41988a <=( a41987a  and  a41984a );
 a41991a <=( (not A298)  and  (not A268) );
 a41994a <=( (not A301)  and  (not A299) );
 a41995a <=( a41994a  and  a41991a );
 a41996a <=( a41995a  and  a41988a );
 a42000a <=( (not A166)  and  (not A167) );
 a42001a <=( (not A169)  and  a42000a );
 a42004a <=( A201  and  A200 );
 a42007a <=( (not A233)  and  (not A232) );
 a42008a <=( a42007a  and  a42004a );
 a42009a <=( a42008a  and  a42001a );
 a42012a <=( (not A265)  and  (not A235) );
 a42015a <=( (not A268)  and  (not A266) );
 a42016a <=( a42015a  and  a42012a );
 a42019a <=( A299  and  A298 );
 a42022a <=( (not A301)  and  (not A300) );
 a42023a <=( a42022a  and  a42019a );
 a42024a <=( a42023a  and  a42016a );
 a42028a <=( (not A166)  and  (not A167) );
 a42029a <=( (not A169)  and  a42028a );
 a42032a <=( A200  and  (not A199) );
 a42035a <=( (not A234)  and  A203 );
 a42036a <=( a42035a  and  a42032a );
 a42037a <=( a42036a  and  a42029a );
 a42040a <=( (not A236)  and  (not A235) );
 a42043a <=( (not A268)  and  (not A267) );
 a42044a <=( a42043a  and  a42040a );
 a42047a <=( (not A300)  and  (not A269) );
 a42050a <=( (not A302)  and  (not A301) );
 a42051a <=( a42050a  and  a42047a );
 a42052a <=( a42051a  and  a42044a );
 a42056a <=( (not A166)  and  (not A167) );
 a42057a <=( (not A169)  and  a42056a );
 a42060a <=( A200  and  (not A199) );
 a42063a <=( (not A234)  and  A203 );
 a42064a <=( a42063a  and  a42060a );
 a42065a <=( a42064a  and  a42057a );
 a42068a <=( (not A236)  and  (not A235) );
 a42071a <=( (not A268)  and  (not A267) );
 a42072a <=( a42071a  and  a42068a );
 a42075a <=( (not A298)  and  (not A269) );
 a42078a <=( (not A301)  and  (not A299) );
 a42079a <=( a42078a  and  a42075a );
 a42080a <=( a42079a  and  a42072a );
 a42084a <=( (not A166)  and  (not A167) );
 a42085a <=( (not A169)  and  a42084a );
 a42088a <=( A200  and  (not A199) );
 a42091a <=( (not A234)  and  A203 );
 a42092a <=( a42091a  and  a42088a );
 a42093a <=( a42092a  and  a42085a );
 a42096a <=( (not A236)  and  (not A235) );
 a42099a <=( (not A266)  and  (not A265) );
 a42100a <=( a42099a  and  a42096a );
 a42103a <=( (not A300)  and  (not A268) );
 a42106a <=( (not A302)  and  (not A301) );
 a42107a <=( a42106a  and  a42103a );
 a42108a <=( a42107a  and  a42100a );
 a42112a <=( (not A166)  and  (not A167) );
 a42113a <=( (not A169)  and  a42112a );
 a42116a <=( A200  and  (not A199) );
 a42119a <=( (not A234)  and  A203 );
 a42120a <=( a42119a  and  a42116a );
 a42121a <=( a42120a  and  a42113a );
 a42124a <=( (not A236)  and  (not A235) );
 a42127a <=( (not A266)  and  (not A265) );
 a42128a <=( a42127a  and  a42124a );
 a42131a <=( (not A298)  and  (not A268) );
 a42134a <=( (not A301)  and  (not A299) );
 a42135a <=( a42134a  and  a42131a );
 a42136a <=( a42135a  and  a42128a );
 a42140a <=( (not A166)  and  (not A167) );
 a42141a <=( (not A169)  and  a42140a );
 a42144a <=( A200  and  (not A199) );
 a42147a <=( (not A232)  and  A203 );
 a42148a <=( a42147a  and  a42144a );
 a42149a <=( a42148a  and  a42141a );
 a42152a <=( (not A235)  and  (not A233) );
 a42155a <=( (not A268)  and  (not A267) );
 a42156a <=( a42155a  and  a42152a );
 a42159a <=( (not A300)  and  (not A269) );
 a42162a <=( (not A302)  and  (not A301) );
 a42163a <=( a42162a  and  a42159a );
 a42164a <=( a42163a  and  a42156a );
 a42168a <=( (not A166)  and  (not A167) );
 a42169a <=( (not A169)  and  a42168a );
 a42172a <=( A200  and  (not A199) );
 a42175a <=( (not A232)  and  A203 );
 a42176a <=( a42175a  and  a42172a );
 a42177a <=( a42176a  and  a42169a );
 a42180a <=( (not A235)  and  (not A233) );
 a42183a <=( (not A268)  and  (not A267) );
 a42184a <=( a42183a  and  a42180a );
 a42187a <=( (not A298)  and  (not A269) );
 a42190a <=( (not A301)  and  (not A299) );
 a42191a <=( a42190a  and  a42187a );
 a42192a <=( a42191a  and  a42184a );
 a42196a <=( (not A166)  and  (not A167) );
 a42197a <=( (not A169)  and  a42196a );
 a42200a <=( A200  and  (not A199) );
 a42203a <=( (not A232)  and  A203 );
 a42204a <=( a42203a  and  a42200a );
 a42205a <=( a42204a  and  a42197a );
 a42208a <=( (not A235)  and  (not A233) );
 a42211a <=( (not A266)  and  (not A265) );
 a42212a <=( a42211a  and  a42208a );
 a42215a <=( (not A300)  and  (not A268) );
 a42218a <=( (not A302)  and  (not A301) );
 a42219a <=( a42218a  and  a42215a );
 a42220a <=( a42219a  and  a42212a );
 a42224a <=( (not A166)  and  (not A167) );
 a42225a <=( (not A169)  and  a42224a );
 a42228a <=( A200  and  (not A199) );
 a42231a <=( (not A232)  and  A203 );
 a42232a <=( a42231a  and  a42228a );
 a42233a <=( a42232a  and  a42225a );
 a42236a <=( (not A235)  and  (not A233) );
 a42239a <=( (not A266)  and  (not A265) );
 a42240a <=( a42239a  and  a42236a );
 a42243a <=( (not A298)  and  (not A268) );
 a42246a <=( (not A301)  and  (not A299) );
 a42247a <=( a42246a  and  a42243a );
 a42248a <=( a42247a  and  a42240a );
 a42252a <=( (not A166)  and  (not A167) );
 a42253a <=( (not A169)  and  a42252a );
 a42256a <=( (not A200)  and  A199 );
 a42259a <=( (not A234)  and  A203 );
 a42260a <=( a42259a  and  a42256a );
 a42261a <=( a42260a  and  a42253a );
 a42264a <=( (not A236)  and  (not A235) );
 a42267a <=( (not A268)  and  (not A267) );
 a42268a <=( a42267a  and  a42264a );
 a42271a <=( (not A300)  and  (not A269) );
 a42274a <=( (not A302)  and  (not A301) );
 a42275a <=( a42274a  and  a42271a );
 a42276a <=( a42275a  and  a42268a );
 a42280a <=( (not A166)  and  (not A167) );
 a42281a <=( (not A169)  and  a42280a );
 a42284a <=( (not A200)  and  A199 );
 a42287a <=( (not A234)  and  A203 );
 a42288a <=( a42287a  and  a42284a );
 a42289a <=( a42288a  and  a42281a );
 a42292a <=( (not A236)  and  (not A235) );
 a42295a <=( (not A268)  and  (not A267) );
 a42296a <=( a42295a  and  a42292a );
 a42299a <=( (not A298)  and  (not A269) );
 a42302a <=( (not A301)  and  (not A299) );
 a42303a <=( a42302a  and  a42299a );
 a42304a <=( a42303a  and  a42296a );
 a42308a <=( (not A166)  and  (not A167) );
 a42309a <=( (not A169)  and  a42308a );
 a42312a <=( (not A200)  and  A199 );
 a42315a <=( (not A234)  and  A203 );
 a42316a <=( a42315a  and  a42312a );
 a42317a <=( a42316a  and  a42309a );
 a42320a <=( (not A236)  and  (not A235) );
 a42323a <=( (not A266)  and  (not A265) );
 a42324a <=( a42323a  and  a42320a );
 a42327a <=( (not A300)  and  (not A268) );
 a42330a <=( (not A302)  and  (not A301) );
 a42331a <=( a42330a  and  a42327a );
 a42332a <=( a42331a  and  a42324a );
 a42336a <=( (not A166)  and  (not A167) );
 a42337a <=( (not A169)  and  a42336a );
 a42340a <=( (not A200)  and  A199 );
 a42343a <=( (not A234)  and  A203 );
 a42344a <=( a42343a  and  a42340a );
 a42345a <=( a42344a  and  a42337a );
 a42348a <=( (not A236)  and  (not A235) );
 a42351a <=( (not A266)  and  (not A265) );
 a42352a <=( a42351a  and  a42348a );
 a42355a <=( (not A298)  and  (not A268) );
 a42358a <=( (not A301)  and  (not A299) );
 a42359a <=( a42358a  and  a42355a );
 a42360a <=( a42359a  and  a42352a );
 a42364a <=( (not A166)  and  (not A167) );
 a42365a <=( (not A169)  and  a42364a );
 a42368a <=( (not A200)  and  A199 );
 a42371a <=( (not A232)  and  A203 );
 a42372a <=( a42371a  and  a42368a );
 a42373a <=( a42372a  and  a42365a );
 a42376a <=( (not A235)  and  (not A233) );
 a42379a <=( (not A268)  and  (not A267) );
 a42380a <=( a42379a  and  a42376a );
 a42383a <=( (not A300)  and  (not A269) );
 a42386a <=( (not A302)  and  (not A301) );
 a42387a <=( a42386a  and  a42383a );
 a42388a <=( a42387a  and  a42380a );
 a42392a <=( (not A166)  and  (not A167) );
 a42393a <=( (not A169)  and  a42392a );
 a42396a <=( (not A200)  and  A199 );
 a42399a <=( (not A232)  and  A203 );
 a42400a <=( a42399a  and  a42396a );
 a42401a <=( a42400a  and  a42393a );
 a42404a <=( (not A235)  and  (not A233) );
 a42407a <=( (not A268)  and  (not A267) );
 a42408a <=( a42407a  and  a42404a );
 a42411a <=( (not A298)  and  (not A269) );
 a42414a <=( (not A301)  and  (not A299) );
 a42415a <=( a42414a  and  a42411a );
 a42416a <=( a42415a  and  a42408a );
 a42420a <=( (not A166)  and  (not A167) );
 a42421a <=( (not A169)  and  a42420a );
 a42424a <=( (not A200)  and  A199 );
 a42427a <=( (not A232)  and  A203 );
 a42428a <=( a42427a  and  a42424a );
 a42429a <=( a42428a  and  a42421a );
 a42432a <=( (not A235)  and  (not A233) );
 a42435a <=( (not A266)  and  (not A265) );
 a42436a <=( a42435a  and  a42432a );
 a42439a <=( (not A300)  and  (not A268) );
 a42442a <=( (not A302)  and  (not A301) );
 a42443a <=( a42442a  and  a42439a );
 a42444a <=( a42443a  and  a42436a );
 a42448a <=( (not A166)  and  (not A167) );
 a42449a <=( (not A169)  and  a42448a );
 a42452a <=( (not A200)  and  A199 );
 a42455a <=( (not A232)  and  A203 );
 a42456a <=( a42455a  and  a42452a );
 a42457a <=( a42456a  and  a42449a );
 a42460a <=( (not A235)  and  (not A233) );
 a42463a <=( (not A266)  and  (not A265) );
 a42464a <=( a42463a  and  a42460a );
 a42467a <=( (not A298)  and  (not A268) );
 a42470a <=( (not A301)  and  (not A299) );
 a42471a <=( a42470a  and  a42467a );
 a42472a <=( a42471a  and  a42464a );
 a42476a <=( A167  and  (not A168) );
 a42477a <=( (not A169)  and  a42476a );
 a42480a <=( A202  and  A166 );
 a42483a <=( (not A235)  and  (not A234) );
 a42484a <=( a42483a  and  a42480a );
 a42485a <=( a42484a  and  a42477a );
 a42488a <=( (not A267)  and  (not A236) );
 a42491a <=( (not A269)  and  (not A268) );
 a42492a <=( a42491a  and  a42488a );
 a42495a <=( A299  and  A298 );
 a42498a <=( (not A301)  and  (not A300) );
 a42499a <=( a42498a  and  a42495a );
 a42500a <=( a42499a  and  a42492a );
 a42504a <=( A167  and  (not A168) );
 a42505a <=( (not A169)  and  a42504a );
 a42508a <=( A202  and  A166 );
 a42511a <=( (not A235)  and  (not A234) );
 a42512a <=( a42511a  and  a42508a );
 a42513a <=( a42512a  and  a42505a );
 a42516a <=( A265  and  (not A236) );
 a42519a <=( (not A267)  and  A266 );
 a42520a <=( a42519a  and  a42516a );
 a42523a <=( (not A300)  and  (not A268) );
 a42526a <=( (not A302)  and  (not A301) );
 a42527a <=( a42526a  and  a42523a );
 a42528a <=( a42527a  and  a42520a );
 a42532a <=( A167  and  (not A168) );
 a42533a <=( (not A169)  and  a42532a );
 a42536a <=( A202  and  A166 );
 a42539a <=( (not A235)  and  (not A234) );
 a42540a <=( a42539a  and  a42536a );
 a42541a <=( a42540a  and  a42533a );
 a42544a <=( A265  and  (not A236) );
 a42547a <=( (not A267)  and  A266 );
 a42548a <=( a42547a  and  a42544a );
 a42551a <=( (not A298)  and  (not A268) );
 a42554a <=( (not A301)  and  (not A299) );
 a42555a <=( a42554a  and  a42551a );
 a42556a <=( a42555a  and  a42548a );
 a42560a <=( A167  and  (not A168) );
 a42561a <=( (not A169)  and  a42560a );
 a42564a <=( A202  and  A166 );
 a42567a <=( (not A235)  and  (not A234) );
 a42568a <=( a42567a  and  a42564a );
 a42569a <=( a42568a  and  a42561a );
 a42572a <=( (not A265)  and  (not A236) );
 a42575a <=( (not A268)  and  (not A266) );
 a42576a <=( a42575a  and  a42572a );
 a42579a <=( A299  and  A298 );
 a42582a <=( (not A301)  and  (not A300) );
 a42583a <=( a42582a  and  a42579a );
 a42584a <=( a42583a  and  a42576a );
 a42588a <=( A167  and  (not A168) );
 a42589a <=( (not A169)  and  a42588a );
 a42592a <=( A202  and  A166 );
 a42595a <=( A233  and  A232 );
 a42596a <=( a42595a  and  a42592a );
 a42597a <=( a42596a  and  a42589a );
 a42600a <=( (not A235)  and  (not A234) );
 a42603a <=( (not A268)  and  (not A267) );
 a42604a <=( a42603a  and  a42600a );
 a42607a <=( (not A300)  and  (not A269) );
 a42610a <=( (not A302)  and  (not A301) );
 a42611a <=( a42610a  and  a42607a );
 a42612a <=( a42611a  and  a42604a );
 a42616a <=( A167  and  (not A168) );
 a42617a <=( (not A169)  and  a42616a );
 a42620a <=( A202  and  A166 );
 a42623a <=( A233  and  A232 );
 a42624a <=( a42623a  and  a42620a );
 a42625a <=( a42624a  and  a42617a );
 a42628a <=( (not A235)  and  (not A234) );
 a42631a <=( (not A268)  and  (not A267) );
 a42632a <=( a42631a  and  a42628a );
 a42635a <=( (not A298)  and  (not A269) );
 a42638a <=( (not A301)  and  (not A299) );
 a42639a <=( a42638a  and  a42635a );
 a42640a <=( a42639a  and  a42632a );
 a42644a <=( A167  and  (not A168) );
 a42645a <=( (not A169)  and  a42644a );
 a42648a <=( A202  and  A166 );
 a42651a <=( A233  and  A232 );
 a42652a <=( a42651a  and  a42648a );
 a42653a <=( a42652a  and  a42645a );
 a42656a <=( (not A235)  and  (not A234) );
 a42659a <=( (not A266)  and  (not A265) );
 a42660a <=( a42659a  and  a42656a );
 a42663a <=( (not A300)  and  (not A268) );
 a42666a <=( (not A302)  and  (not A301) );
 a42667a <=( a42666a  and  a42663a );
 a42668a <=( a42667a  and  a42660a );
 a42672a <=( A167  and  (not A168) );
 a42673a <=( (not A169)  and  a42672a );
 a42676a <=( A202  and  A166 );
 a42679a <=( A233  and  A232 );
 a42680a <=( a42679a  and  a42676a );
 a42681a <=( a42680a  and  a42673a );
 a42684a <=( (not A235)  and  (not A234) );
 a42687a <=( (not A266)  and  (not A265) );
 a42688a <=( a42687a  and  a42684a );
 a42691a <=( (not A298)  and  (not A268) );
 a42694a <=( (not A301)  and  (not A299) );
 a42695a <=( a42694a  and  a42691a );
 a42696a <=( a42695a  and  a42688a );
 a42700a <=( A167  and  (not A168) );
 a42701a <=( (not A169)  and  a42700a );
 a42704a <=( A202  and  A166 );
 a42707a <=( (not A233)  and  (not A232) );
 a42708a <=( a42707a  and  a42704a );
 a42709a <=( a42708a  and  a42701a );
 a42712a <=( (not A267)  and  (not A235) );
 a42715a <=( (not A269)  and  (not A268) );
 a42716a <=( a42715a  and  a42712a );
 a42719a <=( A299  and  A298 );
 a42722a <=( (not A301)  and  (not A300) );
 a42723a <=( a42722a  and  a42719a );
 a42724a <=( a42723a  and  a42716a );
 a42728a <=( A167  and  (not A168) );
 a42729a <=( (not A169)  and  a42728a );
 a42732a <=( A202  and  A166 );
 a42735a <=( (not A233)  and  (not A232) );
 a42736a <=( a42735a  and  a42732a );
 a42737a <=( a42736a  and  a42729a );
 a42740a <=( A265  and  (not A235) );
 a42743a <=( (not A267)  and  A266 );
 a42744a <=( a42743a  and  a42740a );
 a42747a <=( (not A300)  and  (not A268) );
 a42750a <=( (not A302)  and  (not A301) );
 a42751a <=( a42750a  and  a42747a );
 a42752a <=( a42751a  and  a42744a );
 a42756a <=( A167  and  (not A168) );
 a42757a <=( (not A169)  and  a42756a );
 a42760a <=( A202  and  A166 );
 a42763a <=( (not A233)  and  (not A232) );
 a42764a <=( a42763a  and  a42760a );
 a42765a <=( a42764a  and  a42757a );
 a42768a <=( A265  and  (not A235) );
 a42771a <=( (not A267)  and  A266 );
 a42772a <=( a42771a  and  a42768a );
 a42775a <=( (not A298)  and  (not A268) );
 a42778a <=( (not A301)  and  (not A299) );
 a42779a <=( a42778a  and  a42775a );
 a42780a <=( a42779a  and  a42772a );
 a42784a <=( A167  and  (not A168) );
 a42785a <=( (not A169)  and  a42784a );
 a42788a <=( A202  and  A166 );
 a42791a <=( (not A233)  and  (not A232) );
 a42792a <=( a42791a  and  a42788a );
 a42793a <=( a42792a  and  a42785a );
 a42796a <=( (not A265)  and  (not A235) );
 a42799a <=( (not A268)  and  (not A266) );
 a42800a <=( a42799a  and  a42796a );
 a42803a <=( A299  and  A298 );
 a42806a <=( (not A301)  and  (not A300) );
 a42807a <=( a42806a  and  a42803a );
 a42808a <=( a42807a  and  a42800a );
 a42812a <=( A167  and  (not A168) );
 a42813a <=( (not A169)  and  a42812a );
 a42816a <=( A199  and  A166 );
 a42819a <=( (not A234)  and  A201 );
 a42820a <=( a42819a  and  a42816a );
 a42821a <=( a42820a  and  a42813a );
 a42824a <=( (not A236)  and  (not A235) );
 a42827a <=( (not A268)  and  (not A267) );
 a42828a <=( a42827a  and  a42824a );
 a42831a <=( (not A300)  and  (not A269) );
 a42834a <=( (not A302)  and  (not A301) );
 a42835a <=( a42834a  and  a42831a );
 a42836a <=( a42835a  and  a42828a );
 a42840a <=( A167  and  (not A168) );
 a42841a <=( (not A169)  and  a42840a );
 a42844a <=( A199  and  A166 );
 a42847a <=( (not A234)  and  A201 );
 a42848a <=( a42847a  and  a42844a );
 a42849a <=( a42848a  and  a42841a );
 a42852a <=( (not A236)  and  (not A235) );
 a42855a <=( (not A268)  and  (not A267) );
 a42856a <=( a42855a  and  a42852a );
 a42859a <=( (not A298)  and  (not A269) );
 a42862a <=( (not A301)  and  (not A299) );
 a42863a <=( a42862a  and  a42859a );
 a42864a <=( a42863a  and  a42856a );
 a42868a <=( A167  and  (not A168) );
 a42869a <=( (not A169)  and  a42868a );
 a42872a <=( A199  and  A166 );
 a42875a <=( (not A234)  and  A201 );
 a42876a <=( a42875a  and  a42872a );
 a42877a <=( a42876a  and  a42869a );
 a42880a <=( (not A236)  and  (not A235) );
 a42883a <=( (not A266)  and  (not A265) );
 a42884a <=( a42883a  and  a42880a );
 a42887a <=( (not A300)  and  (not A268) );
 a42890a <=( (not A302)  and  (not A301) );
 a42891a <=( a42890a  and  a42887a );
 a42892a <=( a42891a  and  a42884a );
 a42896a <=( A167  and  (not A168) );
 a42897a <=( (not A169)  and  a42896a );
 a42900a <=( A199  and  A166 );
 a42903a <=( (not A234)  and  A201 );
 a42904a <=( a42903a  and  a42900a );
 a42905a <=( a42904a  and  a42897a );
 a42908a <=( (not A236)  and  (not A235) );
 a42911a <=( (not A266)  and  (not A265) );
 a42912a <=( a42911a  and  a42908a );
 a42915a <=( (not A298)  and  (not A268) );
 a42918a <=( (not A301)  and  (not A299) );
 a42919a <=( a42918a  and  a42915a );
 a42920a <=( a42919a  and  a42912a );
 a42924a <=( A167  and  (not A168) );
 a42925a <=( (not A169)  and  a42924a );
 a42928a <=( A199  and  A166 );
 a42931a <=( (not A232)  and  A201 );
 a42932a <=( a42931a  and  a42928a );
 a42933a <=( a42932a  and  a42925a );
 a42936a <=( (not A235)  and  (not A233) );
 a42939a <=( (not A268)  and  (not A267) );
 a42940a <=( a42939a  and  a42936a );
 a42943a <=( (not A300)  and  (not A269) );
 a42946a <=( (not A302)  and  (not A301) );
 a42947a <=( a42946a  and  a42943a );
 a42948a <=( a42947a  and  a42940a );
 a42952a <=( A167  and  (not A168) );
 a42953a <=( (not A169)  and  a42952a );
 a42956a <=( A199  and  A166 );
 a42959a <=( (not A232)  and  A201 );
 a42960a <=( a42959a  and  a42956a );
 a42961a <=( a42960a  and  a42953a );
 a42964a <=( (not A235)  and  (not A233) );
 a42967a <=( (not A268)  and  (not A267) );
 a42968a <=( a42967a  and  a42964a );
 a42971a <=( (not A298)  and  (not A269) );
 a42974a <=( (not A301)  and  (not A299) );
 a42975a <=( a42974a  and  a42971a );
 a42976a <=( a42975a  and  a42968a );
 a42980a <=( A167  and  (not A168) );
 a42981a <=( (not A169)  and  a42980a );
 a42984a <=( A199  and  A166 );
 a42987a <=( (not A232)  and  A201 );
 a42988a <=( a42987a  and  a42984a );
 a42989a <=( a42988a  and  a42981a );
 a42992a <=( (not A235)  and  (not A233) );
 a42995a <=( (not A266)  and  (not A265) );
 a42996a <=( a42995a  and  a42992a );
 a42999a <=( (not A300)  and  (not A268) );
 a43002a <=( (not A302)  and  (not A301) );
 a43003a <=( a43002a  and  a42999a );
 a43004a <=( a43003a  and  a42996a );
 a43008a <=( A167  and  (not A168) );
 a43009a <=( (not A169)  and  a43008a );
 a43012a <=( A199  and  A166 );
 a43015a <=( (not A232)  and  A201 );
 a43016a <=( a43015a  and  a43012a );
 a43017a <=( a43016a  and  a43009a );
 a43020a <=( (not A235)  and  (not A233) );
 a43023a <=( (not A266)  and  (not A265) );
 a43024a <=( a43023a  and  a43020a );
 a43027a <=( (not A298)  and  (not A268) );
 a43030a <=( (not A301)  and  (not A299) );
 a43031a <=( a43030a  and  a43027a );
 a43032a <=( a43031a  and  a43024a );
 a43036a <=( A167  and  (not A168) );
 a43037a <=( (not A169)  and  a43036a );
 a43040a <=( A200  and  A166 );
 a43043a <=( (not A234)  and  A201 );
 a43044a <=( a43043a  and  a43040a );
 a43045a <=( a43044a  and  a43037a );
 a43048a <=( (not A236)  and  (not A235) );
 a43051a <=( (not A268)  and  (not A267) );
 a43052a <=( a43051a  and  a43048a );
 a43055a <=( (not A300)  and  (not A269) );
 a43058a <=( (not A302)  and  (not A301) );
 a43059a <=( a43058a  and  a43055a );
 a43060a <=( a43059a  and  a43052a );
 a43064a <=( A167  and  (not A168) );
 a43065a <=( (not A169)  and  a43064a );
 a43068a <=( A200  and  A166 );
 a43071a <=( (not A234)  and  A201 );
 a43072a <=( a43071a  and  a43068a );
 a43073a <=( a43072a  and  a43065a );
 a43076a <=( (not A236)  and  (not A235) );
 a43079a <=( (not A268)  and  (not A267) );
 a43080a <=( a43079a  and  a43076a );
 a43083a <=( (not A298)  and  (not A269) );
 a43086a <=( (not A301)  and  (not A299) );
 a43087a <=( a43086a  and  a43083a );
 a43088a <=( a43087a  and  a43080a );
 a43092a <=( A167  and  (not A168) );
 a43093a <=( (not A169)  and  a43092a );
 a43096a <=( A200  and  A166 );
 a43099a <=( (not A234)  and  A201 );
 a43100a <=( a43099a  and  a43096a );
 a43101a <=( a43100a  and  a43093a );
 a43104a <=( (not A236)  and  (not A235) );
 a43107a <=( (not A266)  and  (not A265) );
 a43108a <=( a43107a  and  a43104a );
 a43111a <=( (not A300)  and  (not A268) );
 a43114a <=( (not A302)  and  (not A301) );
 a43115a <=( a43114a  and  a43111a );
 a43116a <=( a43115a  and  a43108a );
 a43120a <=( A167  and  (not A168) );
 a43121a <=( (not A169)  and  a43120a );
 a43124a <=( A200  and  A166 );
 a43127a <=( (not A234)  and  A201 );
 a43128a <=( a43127a  and  a43124a );
 a43129a <=( a43128a  and  a43121a );
 a43132a <=( (not A236)  and  (not A235) );
 a43135a <=( (not A266)  and  (not A265) );
 a43136a <=( a43135a  and  a43132a );
 a43139a <=( (not A298)  and  (not A268) );
 a43142a <=( (not A301)  and  (not A299) );
 a43143a <=( a43142a  and  a43139a );
 a43144a <=( a43143a  and  a43136a );
 a43148a <=( A167  and  (not A168) );
 a43149a <=( (not A169)  and  a43148a );
 a43152a <=( A200  and  A166 );
 a43155a <=( (not A232)  and  A201 );
 a43156a <=( a43155a  and  a43152a );
 a43157a <=( a43156a  and  a43149a );
 a43160a <=( (not A235)  and  (not A233) );
 a43163a <=( (not A268)  and  (not A267) );
 a43164a <=( a43163a  and  a43160a );
 a43167a <=( (not A300)  and  (not A269) );
 a43170a <=( (not A302)  and  (not A301) );
 a43171a <=( a43170a  and  a43167a );
 a43172a <=( a43171a  and  a43164a );
 a43176a <=( A167  and  (not A168) );
 a43177a <=( (not A169)  and  a43176a );
 a43180a <=( A200  and  A166 );
 a43183a <=( (not A232)  and  A201 );
 a43184a <=( a43183a  and  a43180a );
 a43185a <=( a43184a  and  a43177a );
 a43188a <=( (not A235)  and  (not A233) );
 a43191a <=( (not A268)  and  (not A267) );
 a43192a <=( a43191a  and  a43188a );
 a43195a <=( (not A298)  and  (not A269) );
 a43198a <=( (not A301)  and  (not A299) );
 a43199a <=( a43198a  and  a43195a );
 a43200a <=( a43199a  and  a43192a );
 a43204a <=( A167  and  (not A168) );
 a43205a <=( (not A169)  and  a43204a );
 a43208a <=( A200  and  A166 );
 a43211a <=( (not A232)  and  A201 );
 a43212a <=( a43211a  and  a43208a );
 a43213a <=( a43212a  and  a43205a );
 a43216a <=( (not A235)  and  (not A233) );
 a43219a <=( (not A266)  and  (not A265) );
 a43220a <=( a43219a  and  a43216a );
 a43223a <=( (not A300)  and  (not A268) );
 a43226a <=( (not A302)  and  (not A301) );
 a43227a <=( a43226a  and  a43223a );
 a43228a <=( a43227a  and  a43220a );
 a43232a <=( A167  and  (not A168) );
 a43233a <=( (not A169)  and  a43232a );
 a43236a <=( A200  and  A166 );
 a43239a <=( (not A232)  and  A201 );
 a43240a <=( a43239a  and  a43236a );
 a43241a <=( a43240a  and  a43233a );
 a43244a <=( (not A235)  and  (not A233) );
 a43247a <=( (not A266)  and  (not A265) );
 a43248a <=( a43247a  and  a43244a );
 a43251a <=( (not A298)  and  (not A268) );
 a43254a <=( (not A301)  and  (not A299) );
 a43255a <=( a43254a  and  a43251a );
 a43256a <=( a43255a  and  a43248a );
 a43260a <=( (not A168)  and  (not A169) );
 a43261a <=( (not A170)  and  a43260a );
 a43264a <=( (not A234)  and  A202 );
 a43267a <=( (not A236)  and  (not A235) );
 a43268a <=( a43267a  and  a43264a );
 a43269a <=( a43268a  and  a43261a );
 a43272a <=( A266  and  A265 );
 a43275a <=( (not A268)  and  (not A267) );
 a43276a <=( a43275a  and  a43272a );
 a43279a <=( A299  and  A298 );
 a43282a <=( (not A301)  and  (not A300) );
 a43283a <=( a43282a  and  a43279a );
 a43284a <=( a43283a  and  a43276a );
 a43288a <=( (not A168)  and  (not A169) );
 a43289a <=( (not A170)  and  a43288a );
 a43292a <=( A232  and  A202 );
 a43295a <=( (not A234)  and  A233 );
 a43296a <=( a43295a  and  a43292a );
 a43297a <=( a43296a  and  a43289a );
 a43300a <=( (not A267)  and  (not A235) );
 a43303a <=( (not A269)  and  (not A268) );
 a43304a <=( a43303a  and  a43300a );
 a43307a <=( A299  and  A298 );
 a43310a <=( (not A301)  and  (not A300) );
 a43311a <=( a43310a  and  a43307a );
 a43312a <=( a43311a  and  a43304a );
 a43316a <=( (not A168)  and  (not A169) );
 a43317a <=( (not A170)  and  a43316a );
 a43320a <=( A232  and  A202 );
 a43323a <=( (not A234)  and  A233 );
 a43324a <=( a43323a  and  a43320a );
 a43325a <=( a43324a  and  a43317a );
 a43328a <=( A265  and  (not A235) );
 a43331a <=( (not A267)  and  A266 );
 a43332a <=( a43331a  and  a43328a );
 a43335a <=( (not A300)  and  (not A268) );
 a43338a <=( (not A302)  and  (not A301) );
 a43339a <=( a43338a  and  a43335a );
 a43340a <=( a43339a  and  a43332a );
 a43344a <=( (not A168)  and  (not A169) );
 a43345a <=( (not A170)  and  a43344a );
 a43348a <=( A232  and  A202 );
 a43351a <=( (not A234)  and  A233 );
 a43352a <=( a43351a  and  a43348a );
 a43353a <=( a43352a  and  a43345a );
 a43356a <=( A265  and  (not A235) );
 a43359a <=( (not A267)  and  A266 );
 a43360a <=( a43359a  and  a43356a );
 a43363a <=( (not A298)  and  (not A268) );
 a43366a <=( (not A301)  and  (not A299) );
 a43367a <=( a43366a  and  a43363a );
 a43368a <=( a43367a  and  a43360a );
 a43372a <=( (not A168)  and  (not A169) );
 a43373a <=( (not A170)  and  a43372a );
 a43376a <=( A232  and  A202 );
 a43379a <=( (not A234)  and  A233 );
 a43380a <=( a43379a  and  a43376a );
 a43381a <=( a43380a  and  a43373a );
 a43384a <=( (not A265)  and  (not A235) );
 a43387a <=( (not A268)  and  (not A266) );
 a43388a <=( a43387a  and  a43384a );
 a43391a <=( A299  and  A298 );
 a43394a <=( (not A301)  and  (not A300) );
 a43395a <=( a43394a  and  a43391a );
 a43396a <=( a43395a  and  a43388a );
 a43400a <=( (not A168)  and  (not A169) );
 a43401a <=( (not A170)  and  a43400a );
 a43404a <=( (not A232)  and  A202 );
 a43407a <=( (not A235)  and  (not A233) );
 a43408a <=( a43407a  and  a43404a );
 a43409a <=( a43408a  and  a43401a );
 a43412a <=( A266  and  A265 );
 a43415a <=( (not A268)  and  (not A267) );
 a43416a <=( a43415a  and  a43412a );
 a43419a <=( A299  and  A298 );
 a43422a <=( (not A301)  and  (not A300) );
 a43423a <=( a43422a  and  a43419a );
 a43424a <=( a43423a  and  a43416a );
 a43428a <=( (not A168)  and  (not A169) );
 a43429a <=( (not A170)  and  a43428a );
 a43432a <=( A201  and  A199 );
 a43435a <=( (not A235)  and  (not A234) );
 a43436a <=( a43435a  and  a43432a );
 a43437a <=( a43436a  and  a43429a );
 a43440a <=( (not A267)  and  (not A236) );
 a43443a <=( (not A269)  and  (not A268) );
 a43444a <=( a43443a  and  a43440a );
 a43447a <=( A299  and  A298 );
 a43450a <=( (not A301)  and  (not A300) );
 a43451a <=( a43450a  and  a43447a );
 a43452a <=( a43451a  and  a43444a );
 a43456a <=( (not A168)  and  (not A169) );
 a43457a <=( (not A170)  and  a43456a );
 a43460a <=( A201  and  A199 );
 a43463a <=( (not A235)  and  (not A234) );
 a43464a <=( a43463a  and  a43460a );
 a43465a <=( a43464a  and  a43457a );
 a43468a <=( A265  and  (not A236) );
 a43471a <=( (not A267)  and  A266 );
 a43472a <=( a43471a  and  a43468a );
 a43475a <=( (not A300)  and  (not A268) );
 a43478a <=( (not A302)  and  (not A301) );
 a43479a <=( a43478a  and  a43475a );
 a43480a <=( a43479a  and  a43472a );
 a43484a <=( (not A168)  and  (not A169) );
 a43485a <=( (not A170)  and  a43484a );
 a43488a <=( A201  and  A199 );
 a43491a <=( (not A235)  and  (not A234) );
 a43492a <=( a43491a  and  a43488a );
 a43493a <=( a43492a  and  a43485a );
 a43496a <=( A265  and  (not A236) );
 a43499a <=( (not A267)  and  A266 );
 a43500a <=( a43499a  and  a43496a );
 a43503a <=( (not A298)  and  (not A268) );
 a43506a <=( (not A301)  and  (not A299) );
 a43507a <=( a43506a  and  a43503a );
 a43508a <=( a43507a  and  a43500a );
 a43512a <=( (not A168)  and  (not A169) );
 a43513a <=( (not A170)  and  a43512a );
 a43516a <=( A201  and  A199 );
 a43519a <=( (not A235)  and  (not A234) );
 a43520a <=( a43519a  and  a43516a );
 a43521a <=( a43520a  and  a43513a );
 a43524a <=( (not A265)  and  (not A236) );
 a43527a <=( (not A268)  and  (not A266) );
 a43528a <=( a43527a  and  a43524a );
 a43531a <=( A299  and  A298 );
 a43534a <=( (not A301)  and  (not A300) );
 a43535a <=( a43534a  and  a43531a );
 a43536a <=( a43535a  and  a43528a );
 a43540a <=( (not A168)  and  (not A169) );
 a43541a <=( (not A170)  and  a43540a );
 a43544a <=( A201  and  A199 );
 a43547a <=( A233  and  A232 );
 a43548a <=( a43547a  and  a43544a );
 a43549a <=( a43548a  and  a43541a );
 a43552a <=( (not A235)  and  (not A234) );
 a43555a <=( (not A268)  and  (not A267) );
 a43556a <=( a43555a  and  a43552a );
 a43559a <=( (not A300)  and  (not A269) );
 a43562a <=( (not A302)  and  (not A301) );
 a43563a <=( a43562a  and  a43559a );
 a43564a <=( a43563a  and  a43556a );
 a43568a <=( (not A168)  and  (not A169) );
 a43569a <=( (not A170)  and  a43568a );
 a43572a <=( A201  and  A199 );
 a43575a <=( A233  and  A232 );
 a43576a <=( a43575a  and  a43572a );
 a43577a <=( a43576a  and  a43569a );
 a43580a <=( (not A235)  and  (not A234) );
 a43583a <=( (not A268)  and  (not A267) );
 a43584a <=( a43583a  and  a43580a );
 a43587a <=( (not A298)  and  (not A269) );
 a43590a <=( (not A301)  and  (not A299) );
 a43591a <=( a43590a  and  a43587a );
 a43592a <=( a43591a  and  a43584a );
 a43596a <=( (not A168)  and  (not A169) );
 a43597a <=( (not A170)  and  a43596a );
 a43600a <=( A201  and  A199 );
 a43603a <=( A233  and  A232 );
 a43604a <=( a43603a  and  a43600a );
 a43605a <=( a43604a  and  a43597a );
 a43608a <=( (not A235)  and  (not A234) );
 a43611a <=( (not A266)  and  (not A265) );
 a43612a <=( a43611a  and  a43608a );
 a43615a <=( (not A300)  and  (not A268) );
 a43618a <=( (not A302)  and  (not A301) );
 a43619a <=( a43618a  and  a43615a );
 a43620a <=( a43619a  and  a43612a );
 a43624a <=( (not A168)  and  (not A169) );
 a43625a <=( (not A170)  and  a43624a );
 a43628a <=( A201  and  A199 );
 a43631a <=( A233  and  A232 );
 a43632a <=( a43631a  and  a43628a );
 a43633a <=( a43632a  and  a43625a );
 a43636a <=( (not A235)  and  (not A234) );
 a43639a <=( (not A266)  and  (not A265) );
 a43640a <=( a43639a  and  a43636a );
 a43643a <=( (not A298)  and  (not A268) );
 a43646a <=( (not A301)  and  (not A299) );
 a43647a <=( a43646a  and  a43643a );
 a43648a <=( a43647a  and  a43640a );
 a43652a <=( (not A168)  and  (not A169) );
 a43653a <=( (not A170)  and  a43652a );
 a43656a <=( A201  and  A199 );
 a43659a <=( (not A233)  and  (not A232) );
 a43660a <=( a43659a  and  a43656a );
 a43661a <=( a43660a  and  a43653a );
 a43664a <=( (not A267)  and  (not A235) );
 a43667a <=( (not A269)  and  (not A268) );
 a43668a <=( a43667a  and  a43664a );
 a43671a <=( A299  and  A298 );
 a43674a <=( (not A301)  and  (not A300) );
 a43675a <=( a43674a  and  a43671a );
 a43676a <=( a43675a  and  a43668a );
 a43680a <=( (not A168)  and  (not A169) );
 a43681a <=( (not A170)  and  a43680a );
 a43684a <=( A201  and  A199 );
 a43687a <=( (not A233)  and  (not A232) );
 a43688a <=( a43687a  and  a43684a );
 a43689a <=( a43688a  and  a43681a );
 a43692a <=( A265  and  (not A235) );
 a43695a <=( (not A267)  and  A266 );
 a43696a <=( a43695a  and  a43692a );
 a43699a <=( (not A300)  and  (not A268) );
 a43702a <=( (not A302)  and  (not A301) );
 a43703a <=( a43702a  and  a43699a );
 a43704a <=( a43703a  and  a43696a );
 a43708a <=( (not A168)  and  (not A169) );
 a43709a <=( (not A170)  and  a43708a );
 a43712a <=( A201  and  A199 );
 a43715a <=( (not A233)  and  (not A232) );
 a43716a <=( a43715a  and  a43712a );
 a43717a <=( a43716a  and  a43709a );
 a43720a <=( A265  and  (not A235) );
 a43723a <=( (not A267)  and  A266 );
 a43724a <=( a43723a  and  a43720a );
 a43727a <=( (not A298)  and  (not A268) );
 a43730a <=( (not A301)  and  (not A299) );
 a43731a <=( a43730a  and  a43727a );
 a43732a <=( a43731a  and  a43724a );
 a43736a <=( (not A168)  and  (not A169) );
 a43737a <=( (not A170)  and  a43736a );
 a43740a <=( A201  and  A199 );
 a43743a <=( (not A233)  and  (not A232) );
 a43744a <=( a43743a  and  a43740a );
 a43745a <=( a43744a  and  a43737a );
 a43748a <=( (not A265)  and  (not A235) );
 a43751a <=( (not A268)  and  (not A266) );
 a43752a <=( a43751a  and  a43748a );
 a43755a <=( A299  and  A298 );
 a43758a <=( (not A301)  and  (not A300) );
 a43759a <=( a43758a  and  a43755a );
 a43760a <=( a43759a  and  a43752a );
 a43764a <=( (not A168)  and  (not A169) );
 a43765a <=( (not A170)  and  a43764a );
 a43768a <=( A201  and  A200 );
 a43771a <=( (not A235)  and  (not A234) );
 a43772a <=( a43771a  and  a43768a );
 a43773a <=( a43772a  and  a43765a );
 a43776a <=( (not A267)  and  (not A236) );
 a43779a <=( (not A269)  and  (not A268) );
 a43780a <=( a43779a  and  a43776a );
 a43783a <=( A299  and  A298 );
 a43786a <=( (not A301)  and  (not A300) );
 a43787a <=( a43786a  and  a43783a );
 a43788a <=( a43787a  and  a43780a );
 a43792a <=( (not A168)  and  (not A169) );
 a43793a <=( (not A170)  and  a43792a );
 a43796a <=( A201  and  A200 );
 a43799a <=( (not A235)  and  (not A234) );
 a43800a <=( a43799a  and  a43796a );
 a43801a <=( a43800a  and  a43793a );
 a43804a <=( A265  and  (not A236) );
 a43807a <=( (not A267)  and  A266 );
 a43808a <=( a43807a  and  a43804a );
 a43811a <=( (not A300)  and  (not A268) );
 a43814a <=( (not A302)  and  (not A301) );
 a43815a <=( a43814a  and  a43811a );
 a43816a <=( a43815a  and  a43808a );
 a43820a <=( (not A168)  and  (not A169) );
 a43821a <=( (not A170)  and  a43820a );
 a43824a <=( A201  and  A200 );
 a43827a <=( (not A235)  and  (not A234) );
 a43828a <=( a43827a  and  a43824a );
 a43829a <=( a43828a  and  a43821a );
 a43832a <=( A265  and  (not A236) );
 a43835a <=( (not A267)  and  A266 );
 a43836a <=( a43835a  and  a43832a );
 a43839a <=( (not A298)  and  (not A268) );
 a43842a <=( (not A301)  and  (not A299) );
 a43843a <=( a43842a  and  a43839a );
 a43844a <=( a43843a  and  a43836a );
 a43848a <=( (not A168)  and  (not A169) );
 a43849a <=( (not A170)  and  a43848a );
 a43852a <=( A201  and  A200 );
 a43855a <=( (not A235)  and  (not A234) );
 a43856a <=( a43855a  and  a43852a );
 a43857a <=( a43856a  and  a43849a );
 a43860a <=( (not A265)  and  (not A236) );
 a43863a <=( (not A268)  and  (not A266) );
 a43864a <=( a43863a  and  a43860a );
 a43867a <=( A299  and  A298 );
 a43870a <=( (not A301)  and  (not A300) );
 a43871a <=( a43870a  and  a43867a );
 a43872a <=( a43871a  and  a43864a );
 a43876a <=( (not A168)  and  (not A169) );
 a43877a <=( (not A170)  and  a43876a );
 a43880a <=( A201  and  A200 );
 a43883a <=( A233  and  A232 );
 a43884a <=( a43883a  and  a43880a );
 a43885a <=( a43884a  and  a43877a );
 a43888a <=( (not A235)  and  (not A234) );
 a43891a <=( (not A268)  and  (not A267) );
 a43892a <=( a43891a  and  a43888a );
 a43895a <=( (not A300)  and  (not A269) );
 a43898a <=( (not A302)  and  (not A301) );
 a43899a <=( a43898a  and  a43895a );
 a43900a <=( a43899a  and  a43892a );
 a43904a <=( (not A168)  and  (not A169) );
 a43905a <=( (not A170)  and  a43904a );
 a43908a <=( A201  and  A200 );
 a43911a <=( A233  and  A232 );
 a43912a <=( a43911a  and  a43908a );
 a43913a <=( a43912a  and  a43905a );
 a43916a <=( (not A235)  and  (not A234) );
 a43919a <=( (not A268)  and  (not A267) );
 a43920a <=( a43919a  and  a43916a );
 a43923a <=( (not A298)  and  (not A269) );
 a43926a <=( (not A301)  and  (not A299) );
 a43927a <=( a43926a  and  a43923a );
 a43928a <=( a43927a  and  a43920a );
 a43932a <=( (not A168)  and  (not A169) );
 a43933a <=( (not A170)  and  a43932a );
 a43936a <=( A201  and  A200 );
 a43939a <=( A233  and  A232 );
 a43940a <=( a43939a  and  a43936a );
 a43941a <=( a43940a  and  a43933a );
 a43944a <=( (not A235)  and  (not A234) );
 a43947a <=( (not A266)  and  (not A265) );
 a43948a <=( a43947a  and  a43944a );
 a43951a <=( (not A300)  and  (not A268) );
 a43954a <=( (not A302)  and  (not A301) );
 a43955a <=( a43954a  and  a43951a );
 a43956a <=( a43955a  and  a43948a );
 a43960a <=( (not A168)  and  (not A169) );
 a43961a <=( (not A170)  and  a43960a );
 a43964a <=( A201  and  A200 );
 a43967a <=( A233  and  A232 );
 a43968a <=( a43967a  and  a43964a );
 a43969a <=( a43968a  and  a43961a );
 a43972a <=( (not A235)  and  (not A234) );
 a43975a <=( (not A266)  and  (not A265) );
 a43976a <=( a43975a  and  a43972a );
 a43979a <=( (not A298)  and  (not A268) );
 a43982a <=( (not A301)  and  (not A299) );
 a43983a <=( a43982a  and  a43979a );
 a43984a <=( a43983a  and  a43976a );
 a43988a <=( (not A168)  and  (not A169) );
 a43989a <=( (not A170)  and  a43988a );
 a43992a <=( A201  and  A200 );
 a43995a <=( (not A233)  and  (not A232) );
 a43996a <=( a43995a  and  a43992a );
 a43997a <=( a43996a  and  a43989a );
 a44000a <=( (not A267)  and  (not A235) );
 a44003a <=( (not A269)  and  (not A268) );
 a44004a <=( a44003a  and  a44000a );
 a44007a <=( A299  and  A298 );
 a44010a <=( (not A301)  and  (not A300) );
 a44011a <=( a44010a  and  a44007a );
 a44012a <=( a44011a  and  a44004a );
 a44016a <=( (not A168)  and  (not A169) );
 a44017a <=( (not A170)  and  a44016a );
 a44020a <=( A201  and  A200 );
 a44023a <=( (not A233)  and  (not A232) );
 a44024a <=( a44023a  and  a44020a );
 a44025a <=( a44024a  and  a44017a );
 a44028a <=( A265  and  (not A235) );
 a44031a <=( (not A267)  and  A266 );
 a44032a <=( a44031a  and  a44028a );
 a44035a <=( (not A300)  and  (not A268) );
 a44038a <=( (not A302)  and  (not A301) );
 a44039a <=( a44038a  and  a44035a );
 a44040a <=( a44039a  and  a44032a );
 a44044a <=( (not A168)  and  (not A169) );
 a44045a <=( (not A170)  and  a44044a );
 a44048a <=( A201  and  A200 );
 a44051a <=( (not A233)  and  (not A232) );
 a44052a <=( a44051a  and  a44048a );
 a44053a <=( a44052a  and  a44045a );
 a44056a <=( A265  and  (not A235) );
 a44059a <=( (not A267)  and  A266 );
 a44060a <=( a44059a  and  a44056a );
 a44063a <=( (not A298)  and  (not A268) );
 a44066a <=( (not A301)  and  (not A299) );
 a44067a <=( a44066a  and  a44063a );
 a44068a <=( a44067a  and  a44060a );
 a44072a <=( (not A168)  and  (not A169) );
 a44073a <=( (not A170)  and  a44072a );
 a44076a <=( A201  and  A200 );
 a44079a <=( (not A233)  and  (not A232) );
 a44080a <=( a44079a  and  a44076a );
 a44081a <=( a44080a  and  a44073a );
 a44084a <=( (not A265)  and  (not A235) );
 a44087a <=( (not A268)  and  (not A266) );
 a44088a <=( a44087a  and  a44084a );
 a44091a <=( A299  and  A298 );
 a44094a <=( (not A301)  and  (not A300) );
 a44095a <=( a44094a  and  a44091a );
 a44096a <=( a44095a  and  a44088a );
 a44100a <=( (not A168)  and  (not A169) );
 a44101a <=( (not A170)  and  a44100a );
 a44104a <=( A200  and  (not A199) );
 a44107a <=( (not A234)  and  A203 );
 a44108a <=( a44107a  and  a44104a );
 a44109a <=( a44108a  and  a44101a );
 a44112a <=( (not A236)  and  (not A235) );
 a44115a <=( (not A268)  and  (not A267) );
 a44116a <=( a44115a  and  a44112a );
 a44119a <=( (not A300)  and  (not A269) );
 a44122a <=( (not A302)  and  (not A301) );
 a44123a <=( a44122a  and  a44119a );
 a44124a <=( a44123a  and  a44116a );
 a44128a <=( (not A168)  and  (not A169) );
 a44129a <=( (not A170)  and  a44128a );
 a44132a <=( A200  and  (not A199) );
 a44135a <=( (not A234)  and  A203 );
 a44136a <=( a44135a  and  a44132a );
 a44137a <=( a44136a  and  a44129a );
 a44140a <=( (not A236)  and  (not A235) );
 a44143a <=( (not A268)  and  (not A267) );
 a44144a <=( a44143a  and  a44140a );
 a44147a <=( (not A298)  and  (not A269) );
 a44150a <=( (not A301)  and  (not A299) );
 a44151a <=( a44150a  and  a44147a );
 a44152a <=( a44151a  and  a44144a );
 a44156a <=( (not A168)  and  (not A169) );
 a44157a <=( (not A170)  and  a44156a );
 a44160a <=( A200  and  (not A199) );
 a44163a <=( (not A234)  and  A203 );
 a44164a <=( a44163a  and  a44160a );
 a44165a <=( a44164a  and  a44157a );
 a44168a <=( (not A236)  and  (not A235) );
 a44171a <=( (not A266)  and  (not A265) );
 a44172a <=( a44171a  and  a44168a );
 a44175a <=( (not A300)  and  (not A268) );
 a44178a <=( (not A302)  and  (not A301) );
 a44179a <=( a44178a  and  a44175a );
 a44180a <=( a44179a  and  a44172a );
 a44184a <=( (not A168)  and  (not A169) );
 a44185a <=( (not A170)  and  a44184a );
 a44188a <=( A200  and  (not A199) );
 a44191a <=( (not A234)  and  A203 );
 a44192a <=( a44191a  and  a44188a );
 a44193a <=( a44192a  and  a44185a );
 a44196a <=( (not A236)  and  (not A235) );
 a44199a <=( (not A266)  and  (not A265) );
 a44200a <=( a44199a  and  a44196a );
 a44203a <=( (not A298)  and  (not A268) );
 a44206a <=( (not A301)  and  (not A299) );
 a44207a <=( a44206a  and  a44203a );
 a44208a <=( a44207a  and  a44200a );
 a44212a <=( (not A168)  and  (not A169) );
 a44213a <=( (not A170)  and  a44212a );
 a44216a <=( A200  and  (not A199) );
 a44219a <=( (not A232)  and  A203 );
 a44220a <=( a44219a  and  a44216a );
 a44221a <=( a44220a  and  a44213a );
 a44224a <=( (not A235)  and  (not A233) );
 a44227a <=( (not A268)  and  (not A267) );
 a44228a <=( a44227a  and  a44224a );
 a44231a <=( (not A300)  and  (not A269) );
 a44234a <=( (not A302)  and  (not A301) );
 a44235a <=( a44234a  and  a44231a );
 a44236a <=( a44235a  and  a44228a );
 a44240a <=( (not A168)  and  (not A169) );
 a44241a <=( (not A170)  and  a44240a );
 a44244a <=( A200  and  (not A199) );
 a44247a <=( (not A232)  and  A203 );
 a44248a <=( a44247a  and  a44244a );
 a44249a <=( a44248a  and  a44241a );
 a44252a <=( (not A235)  and  (not A233) );
 a44255a <=( (not A268)  and  (not A267) );
 a44256a <=( a44255a  and  a44252a );
 a44259a <=( (not A298)  and  (not A269) );
 a44262a <=( (not A301)  and  (not A299) );
 a44263a <=( a44262a  and  a44259a );
 a44264a <=( a44263a  and  a44256a );
 a44268a <=( (not A168)  and  (not A169) );
 a44269a <=( (not A170)  and  a44268a );
 a44272a <=( A200  and  (not A199) );
 a44275a <=( (not A232)  and  A203 );
 a44276a <=( a44275a  and  a44272a );
 a44277a <=( a44276a  and  a44269a );
 a44280a <=( (not A235)  and  (not A233) );
 a44283a <=( (not A266)  and  (not A265) );
 a44284a <=( a44283a  and  a44280a );
 a44287a <=( (not A300)  and  (not A268) );
 a44290a <=( (not A302)  and  (not A301) );
 a44291a <=( a44290a  and  a44287a );
 a44292a <=( a44291a  and  a44284a );
 a44296a <=( (not A168)  and  (not A169) );
 a44297a <=( (not A170)  and  a44296a );
 a44300a <=( A200  and  (not A199) );
 a44303a <=( (not A232)  and  A203 );
 a44304a <=( a44303a  and  a44300a );
 a44305a <=( a44304a  and  a44297a );
 a44308a <=( (not A235)  and  (not A233) );
 a44311a <=( (not A266)  and  (not A265) );
 a44312a <=( a44311a  and  a44308a );
 a44315a <=( (not A298)  and  (not A268) );
 a44318a <=( (not A301)  and  (not A299) );
 a44319a <=( a44318a  and  a44315a );
 a44320a <=( a44319a  and  a44312a );
 a44324a <=( (not A168)  and  (not A169) );
 a44325a <=( (not A170)  and  a44324a );
 a44328a <=( (not A200)  and  A199 );
 a44331a <=( (not A234)  and  A203 );
 a44332a <=( a44331a  and  a44328a );
 a44333a <=( a44332a  and  a44325a );
 a44336a <=( (not A236)  and  (not A235) );
 a44339a <=( (not A268)  and  (not A267) );
 a44340a <=( a44339a  and  a44336a );
 a44343a <=( (not A300)  and  (not A269) );
 a44346a <=( (not A302)  and  (not A301) );
 a44347a <=( a44346a  and  a44343a );
 a44348a <=( a44347a  and  a44340a );
 a44352a <=( (not A168)  and  (not A169) );
 a44353a <=( (not A170)  and  a44352a );
 a44356a <=( (not A200)  and  A199 );
 a44359a <=( (not A234)  and  A203 );
 a44360a <=( a44359a  and  a44356a );
 a44361a <=( a44360a  and  a44353a );
 a44364a <=( (not A236)  and  (not A235) );
 a44367a <=( (not A268)  and  (not A267) );
 a44368a <=( a44367a  and  a44364a );
 a44371a <=( (not A298)  and  (not A269) );
 a44374a <=( (not A301)  and  (not A299) );
 a44375a <=( a44374a  and  a44371a );
 a44376a <=( a44375a  and  a44368a );
 a44380a <=( (not A168)  and  (not A169) );
 a44381a <=( (not A170)  and  a44380a );
 a44384a <=( (not A200)  and  A199 );
 a44387a <=( (not A234)  and  A203 );
 a44388a <=( a44387a  and  a44384a );
 a44389a <=( a44388a  and  a44381a );
 a44392a <=( (not A236)  and  (not A235) );
 a44395a <=( (not A266)  and  (not A265) );
 a44396a <=( a44395a  and  a44392a );
 a44399a <=( (not A300)  and  (not A268) );
 a44402a <=( (not A302)  and  (not A301) );
 a44403a <=( a44402a  and  a44399a );
 a44404a <=( a44403a  and  a44396a );
 a44408a <=( (not A168)  and  (not A169) );
 a44409a <=( (not A170)  and  a44408a );
 a44412a <=( (not A200)  and  A199 );
 a44415a <=( (not A234)  and  A203 );
 a44416a <=( a44415a  and  a44412a );
 a44417a <=( a44416a  and  a44409a );
 a44420a <=( (not A236)  and  (not A235) );
 a44423a <=( (not A266)  and  (not A265) );
 a44424a <=( a44423a  and  a44420a );
 a44427a <=( (not A298)  and  (not A268) );
 a44430a <=( (not A301)  and  (not A299) );
 a44431a <=( a44430a  and  a44427a );
 a44432a <=( a44431a  and  a44424a );
 a44436a <=( (not A168)  and  (not A169) );
 a44437a <=( (not A170)  and  a44436a );
 a44440a <=( (not A200)  and  A199 );
 a44443a <=( (not A232)  and  A203 );
 a44444a <=( a44443a  and  a44440a );
 a44445a <=( a44444a  and  a44437a );
 a44448a <=( (not A235)  and  (not A233) );
 a44451a <=( (not A268)  and  (not A267) );
 a44452a <=( a44451a  and  a44448a );
 a44455a <=( (not A300)  and  (not A269) );
 a44458a <=( (not A302)  and  (not A301) );
 a44459a <=( a44458a  and  a44455a );
 a44460a <=( a44459a  and  a44452a );
 a44464a <=( (not A168)  and  (not A169) );
 a44465a <=( (not A170)  and  a44464a );
 a44468a <=( (not A200)  and  A199 );
 a44471a <=( (not A232)  and  A203 );
 a44472a <=( a44471a  and  a44468a );
 a44473a <=( a44472a  and  a44465a );
 a44476a <=( (not A235)  and  (not A233) );
 a44479a <=( (not A268)  and  (not A267) );
 a44480a <=( a44479a  and  a44476a );
 a44483a <=( (not A298)  and  (not A269) );
 a44486a <=( (not A301)  and  (not A299) );
 a44487a <=( a44486a  and  a44483a );
 a44488a <=( a44487a  and  a44480a );
 a44492a <=( (not A168)  and  (not A169) );
 a44493a <=( (not A170)  and  a44492a );
 a44496a <=( (not A200)  and  A199 );
 a44499a <=( (not A232)  and  A203 );
 a44500a <=( a44499a  and  a44496a );
 a44501a <=( a44500a  and  a44493a );
 a44504a <=( (not A235)  and  (not A233) );
 a44507a <=( (not A266)  and  (not A265) );
 a44508a <=( a44507a  and  a44504a );
 a44511a <=( (not A300)  and  (not A268) );
 a44514a <=( (not A302)  and  (not A301) );
 a44515a <=( a44514a  and  a44511a );
 a44516a <=( a44515a  and  a44508a );
 a44520a <=( (not A168)  and  (not A169) );
 a44521a <=( (not A170)  and  a44520a );
 a44524a <=( (not A200)  and  A199 );
 a44527a <=( (not A232)  and  A203 );
 a44528a <=( a44527a  and  a44524a );
 a44529a <=( a44528a  and  a44521a );
 a44532a <=( (not A235)  and  (not A233) );
 a44535a <=( (not A266)  and  (not A265) );
 a44536a <=( a44535a  and  a44532a );
 a44539a <=( (not A298)  and  (not A268) );
 a44542a <=( (not A301)  and  (not A299) );
 a44543a <=( a44542a  and  a44539a );
 a44544a <=( a44543a  and  a44536a );
 a44547a <=( A166  and  A168 );
 a44550a <=( (not A202)  and  (not A201) );
 a44551a <=( a44550a  and  a44547a );
 a44554a <=( (not A234)  and  (not A203) );
 a44557a <=( (not A236)  and  (not A235) );
 a44558a <=( a44557a  and  a44554a );
 a44559a <=( a44558a  and  a44551a );
 a44562a <=( A266  and  A265 );
 a44565a <=( (not A268)  and  (not A267) );
 a44566a <=( a44565a  and  a44562a );
 a44569a <=( A299  and  A298 );
 a44572a <=( (not A301)  and  (not A300) );
 a44573a <=( a44572a  and  a44569a );
 a44574a <=( a44573a  and  a44566a );
 a44577a <=( A166  and  A168 );
 a44580a <=( (not A202)  and  (not A201) );
 a44581a <=( a44580a  and  a44577a );
 a44584a <=( A232  and  (not A203) );
 a44587a <=( (not A234)  and  A233 );
 a44588a <=( a44587a  and  a44584a );
 a44589a <=( a44588a  and  a44581a );
 a44592a <=( (not A267)  and  (not A235) );
 a44595a <=( (not A269)  and  (not A268) );
 a44596a <=( a44595a  and  a44592a );
 a44599a <=( A299  and  A298 );
 a44602a <=( (not A301)  and  (not A300) );
 a44603a <=( a44602a  and  a44599a );
 a44604a <=( a44603a  and  a44596a );
 a44607a <=( A166  and  A168 );
 a44610a <=( (not A202)  and  (not A201) );
 a44611a <=( a44610a  and  a44607a );
 a44614a <=( A232  and  (not A203) );
 a44617a <=( (not A234)  and  A233 );
 a44618a <=( a44617a  and  a44614a );
 a44619a <=( a44618a  and  a44611a );
 a44622a <=( A265  and  (not A235) );
 a44625a <=( (not A267)  and  A266 );
 a44626a <=( a44625a  and  a44622a );
 a44629a <=( (not A300)  and  (not A268) );
 a44632a <=( (not A302)  and  (not A301) );
 a44633a <=( a44632a  and  a44629a );
 a44634a <=( a44633a  and  a44626a );
 a44637a <=( A166  and  A168 );
 a44640a <=( (not A202)  and  (not A201) );
 a44641a <=( a44640a  and  a44637a );
 a44644a <=( A232  and  (not A203) );
 a44647a <=( (not A234)  and  A233 );
 a44648a <=( a44647a  and  a44644a );
 a44649a <=( a44648a  and  a44641a );
 a44652a <=( A265  and  (not A235) );
 a44655a <=( (not A267)  and  A266 );
 a44656a <=( a44655a  and  a44652a );
 a44659a <=( (not A298)  and  (not A268) );
 a44662a <=( (not A301)  and  (not A299) );
 a44663a <=( a44662a  and  a44659a );
 a44664a <=( a44663a  and  a44656a );
 a44667a <=( A166  and  A168 );
 a44670a <=( (not A202)  and  (not A201) );
 a44671a <=( a44670a  and  a44667a );
 a44674a <=( A232  and  (not A203) );
 a44677a <=( (not A234)  and  A233 );
 a44678a <=( a44677a  and  a44674a );
 a44679a <=( a44678a  and  a44671a );
 a44682a <=( (not A265)  and  (not A235) );
 a44685a <=( (not A268)  and  (not A266) );
 a44686a <=( a44685a  and  a44682a );
 a44689a <=( A299  and  A298 );
 a44692a <=( (not A301)  and  (not A300) );
 a44693a <=( a44692a  and  a44689a );
 a44694a <=( a44693a  and  a44686a );
 a44697a <=( A166  and  A168 );
 a44700a <=( (not A202)  and  (not A201) );
 a44701a <=( a44700a  and  a44697a );
 a44704a <=( (not A232)  and  (not A203) );
 a44707a <=( (not A235)  and  (not A233) );
 a44708a <=( a44707a  and  a44704a );
 a44709a <=( a44708a  and  a44701a );
 a44712a <=( A266  and  A265 );
 a44715a <=( (not A268)  and  (not A267) );
 a44716a <=( a44715a  and  a44712a );
 a44719a <=( A299  and  A298 );
 a44722a <=( (not A301)  and  (not A300) );
 a44723a <=( a44722a  and  a44719a );
 a44724a <=( a44723a  and  a44716a );
 a44727a <=( A166  and  A168 );
 a44730a <=( A200  and  A199 );
 a44731a <=( a44730a  and  a44727a );
 a44734a <=( (not A202)  and  (not A201) );
 a44737a <=( (not A235)  and  (not A234) );
 a44738a <=( a44737a  and  a44734a );
 a44739a <=( a44738a  and  a44731a );
 a44742a <=( (not A267)  and  (not A236) );
 a44745a <=( (not A269)  and  (not A268) );
 a44746a <=( a44745a  and  a44742a );
 a44749a <=( A299  and  A298 );
 a44752a <=( (not A301)  and  (not A300) );
 a44753a <=( a44752a  and  a44749a );
 a44754a <=( a44753a  and  a44746a );
 a44757a <=( A166  and  A168 );
 a44760a <=( A200  and  A199 );
 a44761a <=( a44760a  and  a44757a );
 a44764a <=( (not A202)  and  (not A201) );
 a44767a <=( (not A235)  and  (not A234) );
 a44768a <=( a44767a  and  a44764a );
 a44769a <=( a44768a  and  a44761a );
 a44772a <=( A265  and  (not A236) );
 a44775a <=( (not A267)  and  A266 );
 a44776a <=( a44775a  and  a44772a );
 a44779a <=( (not A300)  and  (not A268) );
 a44782a <=( (not A302)  and  (not A301) );
 a44783a <=( a44782a  and  a44779a );
 a44784a <=( a44783a  and  a44776a );
 a44787a <=( A166  and  A168 );
 a44790a <=( A200  and  A199 );
 a44791a <=( a44790a  and  a44787a );
 a44794a <=( (not A202)  and  (not A201) );
 a44797a <=( (not A235)  and  (not A234) );
 a44798a <=( a44797a  and  a44794a );
 a44799a <=( a44798a  and  a44791a );
 a44802a <=( A265  and  (not A236) );
 a44805a <=( (not A267)  and  A266 );
 a44806a <=( a44805a  and  a44802a );
 a44809a <=( (not A298)  and  (not A268) );
 a44812a <=( (not A301)  and  (not A299) );
 a44813a <=( a44812a  and  a44809a );
 a44814a <=( a44813a  and  a44806a );
 a44817a <=( A166  and  A168 );
 a44820a <=( A200  and  A199 );
 a44821a <=( a44820a  and  a44817a );
 a44824a <=( (not A202)  and  (not A201) );
 a44827a <=( (not A235)  and  (not A234) );
 a44828a <=( a44827a  and  a44824a );
 a44829a <=( a44828a  and  a44821a );
 a44832a <=( (not A265)  and  (not A236) );
 a44835a <=( (not A268)  and  (not A266) );
 a44836a <=( a44835a  and  a44832a );
 a44839a <=( A299  and  A298 );
 a44842a <=( (not A301)  and  (not A300) );
 a44843a <=( a44842a  and  a44839a );
 a44844a <=( a44843a  and  a44836a );
 a44847a <=( A166  and  A168 );
 a44850a <=( A200  and  A199 );
 a44851a <=( a44850a  and  a44847a );
 a44854a <=( (not A202)  and  (not A201) );
 a44857a <=( A233  and  A232 );
 a44858a <=( a44857a  and  a44854a );
 a44859a <=( a44858a  and  a44851a );
 a44862a <=( (not A235)  and  (not A234) );
 a44865a <=( (not A268)  and  (not A267) );
 a44866a <=( a44865a  and  a44862a );
 a44869a <=( (not A300)  and  (not A269) );
 a44872a <=( (not A302)  and  (not A301) );
 a44873a <=( a44872a  and  a44869a );
 a44874a <=( a44873a  and  a44866a );
 a44877a <=( A166  and  A168 );
 a44880a <=( A200  and  A199 );
 a44881a <=( a44880a  and  a44877a );
 a44884a <=( (not A202)  and  (not A201) );
 a44887a <=( A233  and  A232 );
 a44888a <=( a44887a  and  a44884a );
 a44889a <=( a44888a  and  a44881a );
 a44892a <=( (not A235)  and  (not A234) );
 a44895a <=( (not A268)  and  (not A267) );
 a44896a <=( a44895a  and  a44892a );
 a44899a <=( (not A298)  and  (not A269) );
 a44902a <=( (not A301)  and  (not A299) );
 a44903a <=( a44902a  and  a44899a );
 a44904a <=( a44903a  and  a44896a );
 a44907a <=( A166  and  A168 );
 a44910a <=( A200  and  A199 );
 a44911a <=( a44910a  and  a44907a );
 a44914a <=( (not A202)  and  (not A201) );
 a44917a <=( A233  and  A232 );
 a44918a <=( a44917a  and  a44914a );
 a44919a <=( a44918a  and  a44911a );
 a44922a <=( (not A235)  and  (not A234) );
 a44925a <=( (not A266)  and  (not A265) );
 a44926a <=( a44925a  and  a44922a );
 a44929a <=( (not A300)  and  (not A268) );
 a44932a <=( (not A302)  and  (not A301) );
 a44933a <=( a44932a  and  a44929a );
 a44934a <=( a44933a  and  a44926a );
 a44937a <=( A166  and  A168 );
 a44940a <=( A200  and  A199 );
 a44941a <=( a44940a  and  a44937a );
 a44944a <=( (not A202)  and  (not A201) );
 a44947a <=( A233  and  A232 );
 a44948a <=( a44947a  and  a44944a );
 a44949a <=( a44948a  and  a44941a );
 a44952a <=( (not A235)  and  (not A234) );
 a44955a <=( (not A266)  and  (not A265) );
 a44956a <=( a44955a  and  a44952a );
 a44959a <=( (not A298)  and  (not A268) );
 a44962a <=( (not A301)  and  (not A299) );
 a44963a <=( a44962a  and  a44959a );
 a44964a <=( a44963a  and  a44956a );
 a44967a <=( A166  and  A168 );
 a44970a <=( A200  and  A199 );
 a44971a <=( a44970a  and  a44967a );
 a44974a <=( (not A202)  and  (not A201) );
 a44977a <=( (not A233)  and  (not A232) );
 a44978a <=( a44977a  and  a44974a );
 a44979a <=( a44978a  and  a44971a );
 a44982a <=( (not A267)  and  (not A235) );
 a44985a <=( (not A269)  and  (not A268) );
 a44986a <=( a44985a  and  a44982a );
 a44989a <=( A299  and  A298 );
 a44992a <=( (not A301)  and  (not A300) );
 a44993a <=( a44992a  and  a44989a );
 a44994a <=( a44993a  and  a44986a );
 a44997a <=( A166  and  A168 );
 a45000a <=( A200  and  A199 );
 a45001a <=( a45000a  and  a44997a );
 a45004a <=( (not A202)  and  (not A201) );
 a45007a <=( (not A233)  and  (not A232) );
 a45008a <=( a45007a  and  a45004a );
 a45009a <=( a45008a  and  a45001a );
 a45012a <=( A265  and  (not A235) );
 a45015a <=( (not A267)  and  A266 );
 a45016a <=( a45015a  and  a45012a );
 a45019a <=( (not A300)  and  (not A268) );
 a45022a <=( (not A302)  and  (not A301) );
 a45023a <=( a45022a  and  a45019a );
 a45024a <=( a45023a  and  a45016a );
 a45027a <=( A166  and  A168 );
 a45030a <=( A200  and  A199 );
 a45031a <=( a45030a  and  a45027a );
 a45034a <=( (not A202)  and  (not A201) );
 a45037a <=( (not A233)  and  (not A232) );
 a45038a <=( a45037a  and  a45034a );
 a45039a <=( a45038a  and  a45031a );
 a45042a <=( A265  and  (not A235) );
 a45045a <=( (not A267)  and  A266 );
 a45046a <=( a45045a  and  a45042a );
 a45049a <=( (not A298)  and  (not A268) );
 a45052a <=( (not A301)  and  (not A299) );
 a45053a <=( a45052a  and  a45049a );
 a45054a <=( a45053a  and  a45046a );
 a45057a <=( A166  and  A168 );
 a45060a <=( A200  and  A199 );
 a45061a <=( a45060a  and  a45057a );
 a45064a <=( (not A202)  and  (not A201) );
 a45067a <=( (not A233)  and  (not A232) );
 a45068a <=( a45067a  and  a45064a );
 a45069a <=( a45068a  and  a45061a );
 a45072a <=( (not A265)  and  (not A235) );
 a45075a <=( (not A268)  and  (not A266) );
 a45076a <=( a45075a  and  a45072a );
 a45079a <=( A299  and  A298 );
 a45082a <=( (not A301)  and  (not A300) );
 a45083a <=( a45082a  and  a45079a );
 a45084a <=( a45083a  and  a45076a );
 a45087a <=( A166  and  A168 );
 a45090a <=( (not A200)  and  (not A199) );
 a45091a <=( a45090a  and  a45087a );
 a45094a <=( (not A234)  and  (not A202) );
 a45097a <=( (not A236)  and  (not A235) );
 a45098a <=( a45097a  and  a45094a );
 a45099a <=( a45098a  and  a45091a );
 a45102a <=( A266  and  A265 );
 a45105a <=( (not A268)  and  (not A267) );
 a45106a <=( a45105a  and  a45102a );
 a45109a <=( A299  and  A298 );
 a45112a <=( (not A301)  and  (not A300) );
 a45113a <=( a45112a  and  a45109a );
 a45114a <=( a45113a  and  a45106a );
 a45117a <=( A166  and  A168 );
 a45120a <=( (not A200)  and  (not A199) );
 a45121a <=( a45120a  and  a45117a );
 a45124a <=( A232  and  (not A202) );
 a45127a <=( (not A234)  and  A233 );
 a45128a <=( a45127a  and  a45124a );
 a45129a <=( a45128a  and  a45121a );
 a45132a <=( (not A267)  and  (not A235) );
 a45135a <=( (not A269)  and  (not A268) );
 a45136a <=( a45135a  and  a45132a );
 a45139a <=( A299  and  A298 );
 a45142a <=( (not A301)  and  (not A300) );
 a45143a <=( a45142a  and  a45139a );
 a45144a <=( a45143a  and  a45136a );
 a45147a <=( A166  and  A168 );
 a45150a <=( (not A200)  and  (not A199) );
 a45151a <=( a45150a  and  a45147a );
 a45154a <=( A232  and  (not A202) );
 a45157a <=( (not A234)  and  A233 );
 a45158a <=( a45157a  and  a45154a );
 a45159a <=( a45158a  and  a45151a );
 a45162a <=( A265  and  (not A235) );
 a45165a <=( (not A267)  and  A266 );
 a45166a <=( a45165a  and  a45162a );
 a45169a <=( (not A300)  and  (not A268) );
 a45172a <=( (not A302)  and  (not A301) );
 a45173a <=( a45172a  and  a45169a );
 a45174a <=( a45173a  and  a45166a );
 a45177a <=( A166  and  A168 );
 a45180a <=( (not A200)  and  (not A199) );
 a45181a <=( a45180a  and  a45177a );
 a45184a <=( A232  and  (not A202) );
 a45187a <=( (not A234)  and  A233 );
 a45188a <=( a45187a  and  a45184a );
 a45189a <=( a45188a  and  a45181a );
 a45192a <=( A265  and  (not A235) );
 a45195a <=( (not A267)  and  A266 );
 a45196a <=( a45195a  and  a45192a );
 a45199a <=( (not A298)  and  (not A268) );
 a45202a <=( (not A301)  and  (not A299) );
 a45203a <=( a45202a  and  a45199a );
 a45204a <=( a45203a  and  a45196a );
 a45207a <=( A166  and  A168 );
 a45210a <=( (not A200)  and  (not A199) );
 a45211a <=( a45210a  and  a45207a );
 a45214a <=( A232  and  (not A202) );
 a45217a <=( (not A234)  and  A233 );
 a45218a <=( a45217a  and  a45214a );
 a45219a <=( a45218a  and  a45211a );
 a45222a <=( (not A265)  and  (not A235) );
 a45225a <=( (not A268)  and  (not A266) );
 a45226a <=( a45225a  and  a45222a );
 a45229a <=( A299  and  A298 );
 a45232a <=( (not A301)  and  (not A300) );
 a45233a <=( a45232a  and  a45229a );
 a45234a <=( a45233a  and  a45226a );
 a45237a <=( A166  and  A168 );
 a45240a <=( (not A200)  and  (not A199) );
 a45241a <=( a45240a  and  a45237a );
 a45244a <=( (not A232)  and  (not A202) );
 a45247a <=( (not A235)  and  (not A233) );
 a45248a <=( a45247a  and  a45244a );
 a45249a <=( a45248a  and  a45241a );
 a45252a <=( A266  and  A265 );
 a45255a <=( (not A268)  and  (not A267) );
 a45256a <=( a45255a  and  a45252a );
 a45259a <=( A299  and  A298 );
 a45262a <=( (not A301)  and  (not A300) );
 a45263a <=( a45262a  and  a45259a );
 a45264a <=( a45263a  and  a45256a );
 a45267a <=( A167  and  A168 );
 a45270a <=( (not A202)  and  (not A201) );
 a45271a <=( a45270a  and  a45267a );
 a45274a <=( (not A234)  and  (not A203) );
 a45277a <=( (not A236)  and  (not A235) );
 a45278a <=( a45277a  and  a45274a );
 a45279a <=( a45278a  and  a45271a );
 a45282a <=( A266  and  A265 );
 a45285a <=( (not A268)  and  (not A267) );
 a45286a <=( a45285a  and  a45282a );
 a45289a <=( A299  and  A298 );
 a45292a <=( (not A301)  and  (not A300) );
 a45293a <=( a45292a  and  a45289a );
 a45294a <=( a45293a  and  a45286a );
 a45297a <=( A167  and  A168 );
 a45300a <=( (not A202)  and  (not A201) );
 a45301a <=( a45300a  and  a45297a );
 a45304a <=( A232  and  (not A203) );
 a45307a <=( (not A234)  and  A233 );
 a45308a <=( a45307a  and  a45304a );
 a45309a <=( a45308a  and  a45301a );
 a45312a <=( (not A267)  and  (not A235) );
 a45315a <=( (not A269)  and  (not A268) );
 a45316a <=( a45315a  and  a45312a );
 a45319a <=( A299  and  A298 );
 a45322a <=( (not A301)  and  (not A300) );
 a45323a <=( a45322a  and  a45319a );
 a45324a <=( a45323a  and  a45316a );
 a45327a <=( A167  and  A168 );
 a45330a <=( (not A202)  and  (not A201) );
 a45331a <=( a45330a  and  a45327a );
 a45334a <=( A232  and  (not A203) );
 a45337a <=( (not A234)  and  A233 );
 a45338a <=( a45337a  and  a45334a );
 a45339a <=( a45338a  and  a45331a );
 a45342a <=( A265  and  (not A235) );
 a45345a <=( (not A267)  and  A266 );
 a45346a <=( a45345a  and  a45342a );
 a45349a <=( (not A300)  and  (not A268) );
 a45352a <=( (not A302)  and  (not A301) );
 a45353a <=( a45352a  and  a45349a );
 a45354a <=( a45353a  and  a45346a );
 a45357a <=( A167  and  A168 );
 a45360a <=( (not A202)  and  (not A201) );
 a45361a <=( a45360a  and  a45357a );
 a45364a <=( A232  and  (not A203) );
 a45367a <=( (not A234)  and  A233 );
 a45368a <=( a45367a  and  a45364a );
 a45369a <=( a45368a  and  a45361a );
 a45372a <=( A265  and  (not A235) );
 a45375a <=( (not A267)  and  A266 );
 a45376a <=( a45375a  and  a45372a );
 a45379a <=( (not A298)  and  (not A268) );
 a45382a <=( (not A301)  and  (not A299) );
 a45383a <=( a45382a  and  a45379a );
 a45384a <=( a45383a  and  a45376a );
 a45387a <=( A167  and  A168 );
 a45390a <=( (not A202)  and  (not A201) );
 a45391a <=( a45390a  and  a45387a );
 a45394a <=( A232  and  (not A203) );
 a45397a <=( (not A234)  and  A233 );
 a45398a <=( a45397a  and  a45394a );
 a45399a <=( a45398a  and  a45391a );
 a45402a <=( (not A265)  and  (not A235) );
 a45405a <=( (not A268)  and  (not A266) );
 a45406a <=( a45405a  and  a45402a );
 a45409a <=( A299  and  A298 );
 a45412a <=( (not A301)  and  (not A300) );
 a45413a <=( a45412a  and  a45409a );
 a45414a <=( a45413a  and  a45406a );
 a45417a <=( A167  and  A168 );
 a45420a <=( (not A202)  and  (not A201) );
 a45421a <=( a45420a  and  a45417a );
 a45424a <=( (not A232)  and  (not A203) );
 a45427a <=( (not A235)  and  (not A233) );
 a45428a <=( a45427a  and  a45424a );
 a45429a <=( a45428a  and  a45421a );
 a45432a <=( A266  and  A265 );
 a45435a <=( (not A268)  and  (not A267) );
 a45436a <=( a45435a  and  a45432a );
 a45439a <=( A299  and  A298 );
 a45442a <=( (not A301)  and  (not A300) );
 a45443a <=( a45442a  and  a45439a );
 a45444a <=( a45443a  and  a45436a );
 a45447a <=( A167  and  A168 );
 a45450a <=( A200  and  A199 );
 a45451a <=( a45450a  and  a45447a );
 a45454a <=( (not A202)  and  (not A201) );
 a45457a <=( (not A235)  and  (not A234) );
 a45458a <=( a45457a  and  a45454a );
 a45459a <=( a45458a  and  a45451a );
 a45462a <=( (not A267)  and  (not A236) );
 a45465a <=( (not A269)  and  (not A268) );
 a45466a <=( a45465a  and  a45462a );
 a45469a <=( A299  and  A298 );
 a45472a <=( (not A301)  and  (not A300) );
 a45473a <=( a45472a  and  a45469a );
 a45474a <=( a45473a  and  a45466a );
 a45477a <=( A167  and  A168 );
 a45480a <=( A200  and  A199 );
 a45481a <=( a45480a  and  a45477a );
 a45484a <=( (not A202)  and  (not A201) );
 a45487a <=( (not A235)  and  (not A234) );
 a45488a <=( a45487a  and  a45484a );
 a45489a <=( a45488a  and  a45481a );
 a45492a <=( A265  and  (not A236) );
 a45495a <=( (not A267)  and  A266 );
 a45496a <=( a45495a  and  a45492a );
 a45499a <=( (not A300)  and  (not A268) );
 a45502a <=( (not A302)  and  (not A301) );
 a45503a <=( a45502a  and  a45499a );
 a45504a <=( a45503a  and  a45496a );
 a45507a <=( A167  and  A168 );
 a45510a <=( A200  and  A199 );
 a45511a <=( a45510a  and  a45507a );
 a45514a <=( (not A202)  and  (not A201) );
 a45517a <=( (not A235)  and  (not A234) );
 a45518a <=( a45517a  and  a45514a );
 a45519a <=( a45518a  and  a45511a );
 a45522a <=( A265  and  (not A236) );
 a45525a <=( (not A267)  and  A266 );
 a45526a <=( a45525a  and  a45522a );
 a45529a <=( (not A298)  and  (not A268) );
 a45532a <=( (not A301)  and  (not A299) );
 a45533a <=( a45532a  and  a45529a );
 a45534a <=( a45533a  and  a45526a );
 a45537a <=( A167  and  A168 );
 a45540a <=( A200  and  A199 );
 a45541a <=( a45540a  and  a45537a );
 a45544a <=( (not A202)  and  (not A201) );
 a45547a <=( (not A235)  and  (not A234) );
 a45548a <=( a45547a  and  a45544a );
 a45549a <=( a45548a  and  a45541a );
 a45552a <=( (not A265)  and  (not A236) );
 a45555a <=( (not A268)  and  (not A266) );
 a45556a <=( a45555a  and  a45552a );
 a45559a <=( A299  and  A298 );
 a45562a <=( (not A301)  and  (not A300) );
 a45563a <=( a45562a  and  a45559a );
 a45564a <=( a45563a  and  a45556a );
 a45567a <=( A167  and  A168 );
 a45570a <=( A200  and  A199 );
 a45571a <=( a45570a  and  a45567a );
 a45574a <=( (not A202)  and  (not A201) );
 a45577a <=( A233  and  A232 );
 a45578a <=( a45577a  and  a45574a );
 a45579a <=( a45578a  and  a45571a );
 a45582a <=( (not A235)  and  (not A234) );
 a45585a <=( (not A268)  and  (not A267) );
 a45586a <=( a45585a  and  a45582a );
 a45589a <=( (not A300)  and  (not A269) );
 a45592a <=( (not A302)  and  (not A301) );
 a45593a <=( a45592a  and  a45589a );
 a45594a <=( a45593a  and  a45586a );
 a45597a <=( A167  and  A168 );
 a45600a <=( A200  and  A199 );
 a45601a <=( a45600a  and  a45597a );
 a45604a <=( (not A202)  and  (not A201) );
 a45607a <=( A233  and  A232 );
 a45608a <=( a45607a  and  a45604a );
 a45609a <=( a45608a  and  a45601a );
 a45612a <=( (not A235)  and  (not A234) );
 a45615a <=( (not A268)  and  (not A267) );
 a45616a <=( a45615a  and  a45612a );
 a45619a <=( (not A298)  and  (not A269) );
 a45622a <=( (not A301)  and  (not A299) );
 a45623a <=( a45622a  and  a45619a );
 a45624a <=( a45623a  and  a45616a );
 a45627a <=( A167  and  A168 );
 a45630a <=( A200  and  A199 );
 a45631a <=( a45630a  and  a45627a );
 a45634a <=( (not A202)  and  (not A201) );
 a45637a <=( A233  and  A232 );
 a45638a <=( a45637a  and  a45634a );
 a45639a <=( a45638a  and  a45631a );
 a45642a <=( (not A235)  and  (not A234) );
 a45645a <=( (not A266)  and  (not A265) );
 a45646a <=( a45645a  and  a45642a );
 a45649a <=( (not A300)  and  (not A268) );
 a45652a <=( (not A302)  and  (not A301) );
 a45653a <=( a45652a  and  a45649a );
 a45654a <=( a45653a  and  a45646a );
 a45657a <=( A167  and  A168 );
 a45660a <=( A200  and  A199 );
 a45661a <=( a45660a  and  a45657a );
 a45664a <=( (not A202)  and  (not A201) );
 a45667a <=( A233  and  A232 );
 a45668a <=( a45667a  and  a45664a );
 a45669a <=( a45668a  and  a45661a );
 a45672a <=( (not A235)  and  (not A234) );
 a45675a <=( (not A266)  and  (not A265) );
 a45676a <=( a45675a  and  a45672a );
 a45679a <=( (not A298)  and  (not A268) );
 a45682a <=( (not A301)  and  (not A299) );
 a45683a <=( a45682a  and  a45679a );
 a45684a <=( a45683a  and  a45676a );
 a45687a <=( A167  and  A168 );
 a45690a <=( A200  and  A199 );
 a45691a <=( a45690a  and  a45687a );
 a45694a <=( (not A202)  and  (not A201) );
 a45697a <=( (not A233)  and  (not A232) );
 a45698a <=( a45697a  and  a45694a );
 a45699a <=( a45698a  and  a45691a );
 a45702a <=( (not A267)  and  (not A235) );
 a45705a <=( (not A269)  and  (not A268) );
 a45706a <=( a45705a  and  a45702a );
 a45709a <=( A299  and  A298 );
 a45712a <=( (not A301)  and  (not A300) );
 a45713a <=( a45712a  and  a45709a );
 a45714a <=( a45713a  and  a45706a );
 a45717a <=( A167  and  A168 );
 a45720a <=( A200  and  A199 );
 a45721a <=( a45720a  and  a45717a );
 a45724a <=( (not A202)  and  (not A201) );
 a45727a <=( (not A233)  and  (not A232) );
 a45728a <=( a45727a  and  a45724a );
 a45729a <=( a45728a  and  a45721a );
 a45732a <=( A265  and  (not A235) );
 a45735a <=( (not A267)  and  A266 );
 a45736a <=( a45735a  and  a45732a );
 a45739a <=( (not A300)  and  (not A268) );
 a45742a <=( (not A302)  and  (not A301) );
 a45743a <=( a45742a  and  a45739a );
 a45744a <=( a45743a  and  a45736a );
 a45747a <=( A167  and  A168 );
 a45750a <=( A200  and  A199 );
 a45751a <=( a45750a  and  a45747a );
 a45754a <=( (not A202)  and  (not A201) );
 a45757a <=( (not A233)  and  (not A232) );
 a45758a <=( a45757a  and  a45754a );
 a45759a <=( a45758a  and  a45751a );
 a45762a <=( A265  and  (not A235) );
 a45765a <=( (not A267)  and  A266 );
 a45766a <=( a45765a  and  a45762a );
 a45769a <=( (not A298)  and  (not A268) );
 a45772a <=( (not A301)  and  (not A299) );
 a45773a <=( a45772a  and  a45769a );
 a45774a <=( a45773a  and  a45766a );
 a45777a <=( A167  and  A168 );
 a45780a <=( A200  and  A199 );
 a45781a <=( a45780a  and  a45777a );
 a45784a <=( (not A202)  and  (not A201) );
 a45787a <=( (not A233)  and  (not A232) );
 a45788a <=( a45787a  and  a45784a );
 a45789a <=( a45788a  and  a45781a );
 a45792a <=( (not A265)  and  (not A235) );
 a45795a <=( (not A268)  and  (not A266) );
 a45796a <=( a45795a  and  a45792a );
 a45799a <=( A299  and  A298 );
 a45802a <=( (not A301)  and  (not A300) );
 a45803a <=( a45802a  and  a45799a );
 a45804a <=( a45803a  and  a45796a );
 a45807a <=( A167  and  A168 );
 a45810a <=( (not A200)  and  (not A199) );
 a45811a <=( a45810a  and  a45807a );
 a45814a <=( (not A234)  and  (not A202) );
 a45817a <=( (not A236)  and  (not A235) );
 a45818a <=( a45817a  and  a45814a );
 a45819a <=( a45818a  and  a45811a );
 a45822a <=( A266  and  A265 );
 a45825a <=( (not A268)  and  (not A267) );
 a45826a <=( a45825a  and  a45822a );
 a45829a <=( A299  and  A298 );
 a45832a <=( (not A301)  and  (not A300) );
 a45833a <=( a45832a  and  a45829a );
 a45834a <=( a45833a  and  a45826a );
 a45837a <=( A167  and  A168 );
 a45840a <=( (not A200)  and  (not A199) );
 a45841a <=( a45840a  and  a45837a );
 a45844a <=( A232  and  (not A202) );
 a45847a <=( (not A234)  and  A233 );
 a45848a <=( a45847a  and  a45844a );
 a45849a <=( a45848a  and  a45841a );
 a45852a <=( (not A267)  and  (not A235) );
 a45855a <=( (not A269)  and  (not A268) );
 a45856a <=( a45855a  and  a45852a );
 a45859a <=( A299  and  A298 );
 a45862a <=( (not A301)  and  (not A300) );
 a45863a <=( a45862a  and  a45859a );
 a45864a <=( a45863a  and  a45856a );
 a45867a <=( A167  and  A168 );
 a45870a <=( (not A200)  and  (not A199) );
 a45871a <=( a45870a  and  a45867a );
 a45874a <=( A232  and  (not A202) );
 a45877a <=( (not A234)  and  A233 );
 a45878a <=( a45877a  and  a45874a );
 a45879a <=( a45878a  and  a45871a );
 a45882a <=( A265  and  (not A235) );
 a45885a <=( (not A267)  and  A266 );
 a45886a <=( a45885a  and  a45882a );
 a45889a <=( (not A300)  and  (not A268) );
 a45892a <=( (not A302)  and  (not A301) );
 a45893a <=( a45892a  and  a45889a );
 a45894a <=( a45893a  and  a45886a );
 a45897a <=( A167  and  A168 );
 a45900a <=( (not A200)  and  (not A199) );
 a45901a <=( a45900a  and  a45897a );
 a45904a <=( A232  and  (not A202) );
 a45907a <=( (not A234)  and  A233 );
 a45908a <=( a45907a  and  a45904a );
 a45909a <=( a45908a  and  a45901a );
 a45912a <=( A265  and  (not A235) );
 a45915a <=( (not A267)  and  A266 );
 a45916a <=( a45915a  and  a45912a );
 a45919a <=( (not A298)  and  (not A268) );
 a45922a <=( (not A301)  and  (not A299) );
 a45923a <=( a45922a  and  a45919a );
 a45924a <=( a45923a  and  a45916a );
 a45927a <=( A167  and  A168 );
 a45930a <=( (not A200)  and  (not A199) );
 a45931a <=( a45930a  and  a45927a );
 a45934a <=( A232  and  (not A202) );
 a45937a <=( (not A234)  and  A233 );
 a45938a <=( a45937a  and  a45934a );
 a45939a <=( a45938a  and  a45931a );
 a45942a <=( (not A265)  and  (not A235) );
 a45945a <=( (not A268)  and  (not A266) );
 a45946a <=( a45945a  and  a45942a );
 a45949a <=( A299  and  A298 );
 a45952a <=( (not A301)  and  (not A300) );
 a45953a <=( a45952a  and  a45949a );
 a45954a <=( a45953a  and  a45946a );
 a45957a <=( A167  and  A168 );
 a45960a <=( (not A200)  and  (not A199) );
 a45961a <=( a45960a  and  a45957a );
 a45964a <=( (not A232)  and  (not A202) );
 a45967a <=( (not A235)  and  (not A233) );
 a45968a <=( a45967a  and  a45964a );
 a45969a <=( a45968a  and  a45961a );
 a45972a <=( A266  and  A265 );
 a45975a <=( (not A268)  and  (not A267) );
 a45976a <=( a45975a  and  a45972a );
 a45979a <=( A299  and  A298 );
 a45982a <=( (not A301)  and  (not A300) );
 a45983a <=( a45982a  and  a45979a );
 a45984a <=( a45983a  and  a45976a );
 a45987a <=( A167  and  A170 );
 a45990a <=( (not A201)  and  (not A166) );
 a45991a <=( a45990a  and  a45987a );
 a45994a <=( (not A203)  and  (not A202) );
 a45997a <=( (not A235)  and  (not A234) );
 a45998a <=( a45997a  and  a45994a );
 a45999a <=( a45998a  and  a45991a );
 a46002a <=( (not A267)  and  (not A236) );
 a46005a <=( (not A269)  and  (not A268) );
 a46006a <=( a46005a  and  a46002a );
 a46009a <=( A299  and  A298 );
 a46012a <=( (not A301)  and  (not A300) );
 a46013a <=( a46012a  and  a46009a );
 a46014a <=( a46013a  and  a46006a );
 a46017a <=( A167  and  A170 );
 a46020a <=( (not A201)  and  (not A166) );
 a46021a <=( a46020a  and  a46017a );
 a46024a <=( (not A203)  and  (not A202) );
 a46027a <=( (not A235)  and  (not A234) );
 a46028a <=( a46027a  and  a46024a );
 a46029a <=( a46028a  and  a46021a );
 a46032a <=( A265  and  (not A236) );
 a46035a <=( (not A267)  and  A266 );
 a46036a <=( a46035a  and  a46032a );
 a46039a <=( (not A300)  and  (not A268) );
 a46042a <=( (not A302)  and  (not A301) );
 a46043a <=( a46042a  and  a46039a );
 a46044a <=( a46043a  and  a46036a );
 a46047a <=( A167  and  A170 );
 a46050a <=( (not A201)  and  (not A166) );
 a46051a <=( a46050a  and  a46047a );
 a46054a <=( (not A203)  and  (not A202) );
 a46057a <=( (not A235)  and  (not A234) );
 a46058a <=( a46057a  and  a46054a );
 a46059a <=( a46058a  and  a46051a );
 a46062a <=( A265  and  (not A236) );
 a46065a <=( (not A267)  and  A266 );
 a46066a <=( a46065a  and  a46062a );
 a46069a <=( (not A298)  and  (not A268) );
 a46072a <=( (not A301)  and  (not A299) );
 a46073a <=( a46072a  and  a46069a );
 a46074a <=( a46073a  and  a46066a );
 a46077a <=( A167  and  A170 );
 a46080a <=( (not A201)  and  (not A166) );
 a46081a <=( a46080a  and  a46077a );
 a46084a <=( (not A203)  and  (not A202) );
 a46087a <=( (not A235)  and  (not A234) );
 a46088a <=( a46087a  and  a46084a );
 a46089a <=( a46088a  and  a46081a );
 a46092a <=( (not A265)  and  (not A236) );
 a46095a <=( (not A268)  and  (not A266) );
 a46096a <=( a46095a  and  a46092a );
 a46099a <=( A299  and  A298 );
 a46102a <=( (not A301)  and  (not A300) );
 a46103a <=( a46102a  and  a46099a );
 a46104a <=( a46103a  and  a46096a );
 a46107a <=( A167  and  A170 );
 a46110a <=( (not A201)  and  (not A166) );
 a46111a <=( a46110a  and  a46107a );
 a46114a <=( (not A203)  and  (not A202) );
 a46117a <=( A233  and  A232 );
 a46118a <=( a46117a  and  a46114a );
 a46119a <=( a46118a  and  a46111a );
 a46122a <=( (not A235)  and  (not A234) );
 a46125a <=( (not A268)  and  (not A267) );
 a46126a <=( a46125a  and  a46122a );
 a46129a <=( (not A300)  and  (not A269) );
 a46132a <=( (not A302)  and  (not A301) );
 a46133a <=( a46132a  and  a46129a );
 a46134a <=( a46133a  and  a46126a );
 a46137a <=( A167  and  A170 );
 a46140a <=( (not A201)  and  (not A166) );
 a46141a <=( a46140a  and  a46137a );
 a46144a <=( (not A203)  and  (not A202) );
 a46147a <=( A233  and  A232 );
 a46148a <=( a46147a  and  a46144a );
 a46149a <=( a46148a  and  a46141a );
 a46152a <=( (not A235)  and  (not A234) );
 a46155a <=( (not A268)  and  (not A267) );
 a46156a <=( a46155a  and  a46152a );
 a46159a <=( (not A298)  and  (not A269) );
 a46162a <=( (not A301)  and  (not A299) );
 a46163a <=( a46162a  and  a46159a );
 a46164a <=( a46163a  and  a46156a );
 a46167a <=( A167  and  A170 );
 a46170a <=( (not A201)  and  (not A166) );
 a46171a <=( a46170a  and  a46167a );
 a46174a <=( (not A203)  and  (not A202) );
 a46177a <=( A233  and  A232 );
 a46178a <=( a46177a  and  a46174a );
 a46179a <=( a46178a  and  a46171a );
 a46182a <=( (not A235)  and  (not A234) );
 a46185a <=( (not A266)  and  (not A265) );
 a46186a <=( a46185a  and  a46182a );
 a46189a <=( (not A300)  and  (not A268) );
 a46192a <=( (not A302)  and  (not A301) );
 a46193a <=( a46192a  and  a46189a );
 a46194a <=( a46193a  and  a46186a );
 a46197a <=( A167  and  A170 );
 a46200a <=( (not A201)  and  (not A166) );
 a46201a <=( a46200a  and  a46197a );
 a46204a <=( (not A203)  and  (not A202) );
 a46207a <=( A233  and  A232 );
 a46208a <=( a46207a  and  a46204a );
 a46209a <=( a46208a  and  a46201a );
 a46212a <=( (not A235)  and  (not A234) );
 a46215a <=( (not A266)  and  (not A265) );
 a46216a <=( a46215a  and  a46212a );
 a46219a <=( (not A298)  and  (not A268) );
 a46222a <=( (not A301)  and  (not A299) );
 a46223a <=( a46222a  and  a46219a );
 a46224a <=( a46223a  and  a46216a );
 a46227a <=( A167  and  A170 );
 a46230a <=( (not A201)  and  (not A166) );
 a46231a <=( a46230a  and  a46227a );
 a46234a <=( (not A203)  and  (not A202) );
 a46237a <=( (not A233)  and  (not A232) );
 a46238a <=( a46237a  and  a46234a );
 a46239a <=( a46238a  and  a46231a );
 a46242a <=( (not A267)  and  (not A235) );
 a46245a <=( (not A269)  and  (not A268) );
 a46246a <=( a46245a  and  a46242a );
 a46249a <=( A299  and  A298 );
 a46252a <=( (not A301)  and  (not A300) );
 a46253a <=( a46252a  and  a46249a );
 a46254a <=( a46253a  and  a46246a );
 a46257a <=( A167  and  A170 );
 a46260a <=( (not A201)  and  (not A166) );
 a46261a <=( a46260a  and  a46257a );
 a46264a <=( (not A203)  and  (not A202) );
 a46267a <=( (not A233)  and  (not A232) );
 a46268a <=( a46267a  and  a46264a );
 a46269a <=( a46268a  and  a46261a );
 a46272a <=( A265  and  (not A235) );
 a46275a <=( (not A267)  and  A266 );
 a46276a <=( a46275a  and  a46272a );
 a46279a <=( (not A300)  and  (not A268) );
 a46282a <=( (not A302)  and  (not A301) );
 a46283a <=( a46282a  and  a46279a );
 a46284a <=( a46283a  and  a46276a );
 a46287a <=( A167  and  A170 );
 a46290a <=( (not A201)  and  (not A166) );
 a46291a <=( a46290a  and  a46287a );
 a46294a <=( (not A203)  and  (not A202) );
 a46297a <=( (not A233)  and  (not A232) );
 a46298a <=( a46297a  and  a46294a );
 a46299a <=( a46298a  and  a46291a );
 a46302a <=( A265  and  (not A235) );
 a46305a <=( (not A267)  and  A266 );
 a46306a <=( a46305a  and  a46302a );
 a46309a <=( (not A298)  and  (not A268) );
 a46312a <=( (not A301)  and  (not A299) );
 a46313a <=( a46312a  and  a46309a );
 a46314a <=( a46313a  and  a46306a );
 a46317a <=( A167  and  A170 );
 a46320a <=( (not A201)  and  (not A166) );
 a46321a <=( a46320a  and  a46317a );
 a46324a <=( (not A203)  and  (not A202) );
 a46327a <=( (not A233)  and  (not A232) );
 a46328a <=( a46327a  and  a46324a );
 a46329a <=( a46328a  and  a46321a );
 a46332a <=( (not A265)  and  (not A235) );
 a46335a <=( (not A268)  and  (not A266) );
 a46336a <=( a46335a  and  a46332a );
 a46339a <=( A299  and  A298 );
 a46342a <=( (not A301)  and  (not A300) );
 a46343a <=( a46342a  and  a46339a );
 a46344a <=( a46343a  and  a46336a );
 a46347a <=( A167  and  A170 );
 a46350a <=( A199  and  (not A166) );
 a46351a <=( a46350a  and  a46347a );
 a46354a <=( (not A201)  and  A200 );
 a46357a <=( (not A234)  and  (not A202) );
 a46358a <=( a46357a  and  a46354a );
 a46359a <=( a46358a  and  a46351a );
 a46362a <=( (not A236)  and  (not A235) );
 a46365a <=( (not A268)  and  (not A267) );
 a46366a <=( a46365a  and  a46362a );
 a46369a <=( (not A300)  and  (not A269) );
 a46372a <=( (not A302)  and  (not A301) );
 a46373a <=( a46372a  and  a46369a );
 a46374a <=( a46373a  and  a46366a );
 a46377a <=( A167  and  A170 );
 a46380a <=( A199  and  (not A166) );
 a46381a <=( a46380a  and  a46377a );
 a46384a <=( (not A201)  and  A200 );
 a46387a <=( (not A234)  and  (not A202) );
 a46388a <=( a46387a  and  a46384a );
 a46389a <=( a46388a  and  a46381a );
 a46392a <=( (not A236)  and  (not A235) );
 a46395a <=( (not A268)  and  (not A267) );
 a46396a <=( a46395a  and  a46392a );
 a46399a <=( (not A298)  and  (not A269) );
 a46402a <=( (not A301)  and  (not A299) );
 a46403a <=( a46402a  and  a46399a );
 a46404a <=( a46403a  and  a46396a );
 a46407a <=( A167  and  A170 );
 a46410a <=( A199  and  (not A166) );
 a46411a <=( a46410a  and  a46407a );
 a46414a <=( (not A201)  and  A200 );
 a46417a <=( (not A234)  and  (not A202) );
 a46418a <=( a46417a  and  a46414a );
 a46419a <=( a46418a  and  a46411a );
 a46422a <=( (not A236)  and  (not A235) );
 a46425a <=( (not A266)  and  (not A265) );
 a46426a <=( a46425a  and  a46422a );
 a46429a <=( (not A300)  and  (not A268) );
 a46432a <=( (not A302)  and  (not A301) );
 a46433a <=( a46432a  and  a46429a );
 a46434a <=( a46433a  and  a46426a );
 a46437a <=( A167  and  A170 );
 a46440a <=( A199  and  (not A166) );
 a46441a <=( a46440a  and  a46437a );
 a46444a <=( (not A201)  and  A200 );
 a46447a <=( (not A234)  and  (not A202) );
 a46448a <=( a46447a  and  a46444a );
 a46449a <=( a46448a  and  a46441a );
 a46452a <=( (not A236)  and  (not A235) );
 a46455a <=( (not A266)  and  (not A265) );
 a46456a <=( a46455a  and  a46452a );
 a46459a <=( (not A298)  and  (not A268) );
 a46462a <=( (not A301)  and  (not A299) );
 a46463a <=( a46462a  and  a46459a );
 a46464a <=( a46463a  and  a46456a );
 a46467a <=( A167  and  A170 );
 a46470a <=( A199  and  (not A166) );
 a46471a <=( a46470a  and  a46467a );
 a46474a <=( (not A201)  and  A200 );
 a46477a <=( (not A232)  and  (not A202) );
 a46478a <=( a46477a  and  a46474a );
 a46479a <=( a46478a  and  a46471a );
 a46482a <=( (not A235)  and  (not A233) );
 a46485a <=( (not A268)  and  (not A267) );
 a46486a <=( a46485a  and  a46482a );
 a46489a <=( (not A300)  and  (not A269) );
 a46492a <=( (not A302)  and  (not A301) );
 a46493a <=( a46492a  and  a46489a );
 a46494a <=( a46493a  and  a46486a );
 a46497a <=( A167  and  A170 );
 a46500a <=( A199  and  (not A166) );
 a46501a <=( a46500a  and  a46497a );
 a46504a <=( (not A201)  and  A200 );
 a46507a <=( (not A232)  and  (not A202) );
 a46508a <=( a46507a  and  a46504a );
 a46509a <=( a46508a  and  a46501a );
 a46512a <=( (not A235)  and  (not A233) );
 a46515a <=( (not A268)  and  (not A267) );
 a46516a <=( a46515a  and  a46512a );
 a46519a <=( (not A298)  and  (not A269) );
 a46522a <=( (not A301)  and  (not A299) );
 a46523a <=( a46522a  and  a46519a );
 a46524a <=( a46523a  and  a46516a );
 a46527a <=( A167  and  A170 );
 a46530a <=( A199  and  (not A166) );
 a46531a <=( a46530a  and  a46527a );
 a46534a <=( (not A201)  and  A200 );
 a46537a <=( (not A232)  and  (not A202) );
 a46538a <=( a46537a  and  a46534a );
 a46539a <=( a46538a  and  a46531a );
 a46542a <=( (not A235)  and  (not A233) );
 a46545a <=( (not A266)  and  (not A265) );
 a46546a <=( a46545a  and  a46542a );
 a46549a <=( (not A300)  and  (not A268) );
 a46552a <=( (not A302)  and  (not A301) );
 a46553a <=( a46552a  and  a46549a );
 a46554a <=( a46553a  and  a46546a );
 a46557a <=( A167  and  A170 );
 a46560a <=( A199  and  (not A166) );
 a46561a <=( a46560a  and  a46557a );
 a46564a <=( (not A201)  and  A200 );
 a46567a <=( (not A232)  and  (not A202) );
 a46568a <=( a46567a  and  a46564a );
 a46569a <=( a46568a  and  a46561a );
 a46572a <=( (not A235)  and  (not A233) );
 a46575a <=( (not A266)  and  (not A265) );
 a46576a <=( a46575a  and  a46572a );
 a46579a <=( (not A298)  and  (not A268) );
 a46582a <=( (not A301)  and  (not A299) );
 a46583a <=( a46582a  and  a46579a );
 a46584a <=( a46583a  and  a46576a );
 a46587a <=( A167  and  A170 );
 a46590a <=( (not A199)  and  (not A166) );
 a46591a <=( a46590a  and  a46587a );
 a46594a <=( (not A202)  and  (not A200) );
 a46597a <=( (not A235)  and  (not A234) );
 a46598a <=( a46597a  and  a46594a );
 a46599a <=( a46598a  and  a46591a );
 a46602a <=( (not A267)  and  (not A236) );
 a46605a <=( (not A269)  and  (not A268) );
 a46606a <=( a46605a  and  a46602a );
 a46609a <=( A299  and  A298 );
 a46612a <=( (not A301)  and  (not A300) );
 a46613a <=( a46612a  and  a46609a );
 a46614a <=( a46613a  and  a46606a );
 a46617a <=( A167  and  A170 );
 a46620a <=( (not A199)  and  (not A166) );
 a46621a <=( a46620a  and  a46617a );
 a46624a <=( (not A202)  and  (not A200) );
 a46627a <=( (not A235)  and  (not A234) );
 a46628a <=( a46627a  and  a46624a );
 a46629a <=( a46628a  and  a46621a );
 a46632a <=( A265  and  (not A236) );
 a46635a <=( (not A267)  and  A266 );
 a46636a <=( a46635a  and  a46632a );
 a46639a <=( (not A300)  and  (not A268) );
 a46642a <=( (not A302)  and  (not A301) );
 a46643a <=( a46642a  and  a46639a );
 a46644a <=( a46643a  and  a46636a );
 a46647a <=( A167  and  A170 );
 a46650a <=( (not A199)  and  (not A166) );
 a46651a <=( a46650a  and  a46647a );
 a46654a <=( (not A202)  and  (not A200) );
 a46657a <=( (not A235)  and  (not A234) );
 a46658a <=( a46657a  and  a46654a );
 a46659a <=( a46658a  and  a46651a );
 a46662a <=( A265  and  (not A236) );
 a46665a <=( (not A267)  and  A266 );
 a46666a <=( a46665a  and  a46662a );
 a46669a <=( (not A298)  and  (not A268) );
 a46672a <=( (not A301)  and  (not A299) );
 a46673a <=( a46672a  and  a46669a );
 a46674a <=( a46673a  and  a46666a );
 a46677a <=( A167  and  A170 );
 a46680a <=( (not A199)  and  (not A166) );
 a46681a <=( a46680a  and  a46677a );
 a46684a <=( (not A202)  and  (not A200) );
 a46687a <=( (not A235)  and  (not A234) );
 a46688a <=( a46687a  and  a46684a );
 a46689a <=( a46688a  and  a46681a );
 a46692a <=( (not A265)  and  (not A236) );
 a46695a <=( (not A268)  and  (not A266) );
 a46696a <=( a46695a  and  a46692a );
 a46699a <=( A299  and  A298 );
 a46702a <=( (not A301)  and  (not A300) );
 a46703a <=( a46702a  and  a46699a );
 a46704a <=( a46703a  and  a46696a );
 a46707a <=( A167  and  A170 );
 a46710a <=( (not A199)  and  (not A166) );
 a46711a <=( a46710a  and  a46707a );
 a46714a <=( (not A202)  and  (not A200) );
 a46717a <=( A233  and  A232 );
 a46718a <=( a46717a  and  a46714a );
 a46719a <=( a46718a  and  a46711a );
 a46722a <=( (not A235)  and  (not A234) );
 a46725a <=( (not A268)  and  (not A267) );
 a46726a <=( a46725a  and  a46722a );
 a46729a <=( (not A300)  and  (not A269) );
 a46732a <=( (not A302)  and  (not A301) );
 a46733a <=( a46732a  and  a46729a );
 a46734a <=( a46733a  and  a46726a );
 a46737a <=( A167  and  A170 );
 a46740a <=( (not A199)  and  (not A166) );
 a46741a <=( a46740a  and  a46737a );
 a46744a <=( (not A202)  and  (not A200) );
 a46747a <=( A233  and  A232 );
 a46748a <=( a46747a  and  a46744a );
 a46749a <=( a46748a  and  a46741a );
 a46752a <=( (not A235)  and  (not A234) );
 a46755a <=( (not A268)  and  (not A267) );
 a46756a <=( a46755a  and  a46752a );
 a46759a <=( (not A298)  and  (not A269) );
 a46762a <=( (not A301)  and  (not A299) );
 a46763a <=( a46762a  and  a46759a );
 a46764a <=( a46763a  and  a46756a );
 a46767a <=( A167  and  A170 );
 a46770a <=( (not A199)  and  (not A166) );
 a46771a <=( a46770a  and  a46767a );
 a46774a <=( (not A202)  and  (not A200) );
 a46777a <=( A233  and  A232 );
 a46778a <=( a46777a  and  a46774a );
 a46779a <=( a46778a  and  a46771a );
 a46782a <=( (not A235)  and  (not A234) );
 a46785a <=( (not A266)  and  (not A265) );
 a46786a <=( a46785a  and  a46782a );
 a46789a <=( (not A300)  and  (not A268) );
 a46792a <=( (not A302)  and  (not A301) );
 a46793a <=( a46792a  and  a46789a );
 a46794a <=( a46793a  and  a46786a );
 a46797a <=( A167  and  A170 );
 a46800a <=( (not A199)  and  (not A166) );
 a46801a <=( a46800a  and  a46797a );
 a46804a <=( (not A202)  and  (not A200) );
 a46807a <=( A233  and  A232 );
 a46808a <=( a46807a  and  a46804a );
 a46809a <=( a46808a  and  a46801a );
 a46812a <=( (not A235)  and  (not A234) );
 a46815a <=( (not A266)  and  (not A265) );
 a46816a <=( a46815a  and  a46812a );
 a46819a <=( (not A298)  and  (not A268) );
 a46822a <=( (not A301)  and  (not A299) );
 a46823a <=( a46822a  and  a46819a );
 a46824a <=( a46823a  and  a46816a );
 a46827a <=( A167  and  A170 );
 a46830a <=( (not A199)  and  (not A166) );
 a46831a <=( a46830a  and  a46827a );
 a46834a <=( (not A202)  and  (not A200) );
 a46837a <=( (not A233)  and  (not A232) );
 a46838a <=( a46837a  and  a46834a );
 a46839a <=( a46838a  and  a46831a );
 a46842a <=( (not A267)  and  (not A235) );
 a46845a <=( (not A269)  and  (not A268) );
 a46846a <=( a46845a  and  a46842a );
 a46849a <=( A299  and  A298 );
 a46852a <=( (not A301)  and  (not A300) );
 a46853a <=( a46852a  and  a46849a );
 a46854a <=( a46853a  and  a46846a );
 a46857a <=( A167  and  A170 );
 a46860a <=( (not A199)  and  (not A166) );
 a46861a <=( a46860a  and  a46857a );
 a46864a <=( (not A202)  and  (not A200) );
 a46867a <=( (not A233)  and  (not A232) );
 a46868a <=( a46867a  and  a46864a );
 a46869a <=( a46868a  and  a46861a );
 a46872a <=( A265  and  (not A235) );
 a46875a <=( (not A267)  and  A266 );
 a46876a <=( a46875a  and  a46872a );
 a46879a <=( (not A300)  and  (not A268) );
 a46882a <=( (not A302)  and  (not A301) );
 a46883a <=( a46882a  and  a46879a );
 a46884a <=( a46883a  and  a46876a );
 a46887a <=( A167  and  A170 );
 a46890a <=( (not A199)  and  (not A166) );
 a46891a <=( a46890a  and  a46887a );
 a46894a <=( (not A202)  and  (not A200) );
 a46897a <=( (not A233)  and  (not A232) );
 a46898a <=( a46897a  and  a46894a );
 a46899a <=( a46898a  and  a46891a );
 a46902a <=( A265  and  (not A235) );
 a46905a <=( (not A267)  and  A266 );
 a46906a <=( a46905a  and  a46902a );
 a46909a <=( (not A298)  and  (not A268) );
 a46912a <=( (not A301)  and  (not A299) );
 a46913a <=( a46912a  and  a46909a );
 a46914a <=( a46913a  and  a46906a );
 a46917a <=( A167  and  A170 );
 a46920a <=( (not A199)  and  (not A166) );
 a46921a <=( a46920a  and  a46917a );
 a46924a <=( (not A202)  and  (not A200) );
 a46927a <=( (not A233)  and  (not A232) );
 a46928a <=( a46927a  and  a46924a );
 a46929a <=( a46928a  and  a46921a );
 a46932a <=( (not A265)  and  (not A235) );
 a46935a <=( (not A268)  and  (not A266) );
 a46936a <=( a46935a  and  a46932a );
 a46939a <=( A299  and  A298 );
 a46942a <=( (not A301)  and  (not A300) );
 a46943a <=( a46942a  and  a46939a );
 a46944a <=( a46943a  and  a46936a );
 a46947a <=( (not A167)  and  A170 );
 a46950a <=( (not A201)  and  A166 );
 a46951a <=( a46950a  and  a46947a );
 a46954a <=( (not A203)  and  (not A202) );
 a46957a <=( (not A235)  and  (not A234) );
 a46958a <=( a46957a  and  a46954a );
 a46959a <=( a46958a  and  a46951a );
 a46962a <=( (not A267)  and  (not A236) );
 a46965a <=( (not A269)  and  (not A268) );
 a46966a <=( a46965a  and  a46962a );
 a46969a <=( A299  and  A298 );
 a46972a <=( (not A301)  and  (not A300) );
 a46973a <=( a46972a  and  a46969a );
 a46974a <=( a46973a  and  a46966a );
 a46977a <=( (not A167)  and  A170 );
 a46980a <=( (not A201)  and  A166 );
 a46981a <=( a46980a  and  a46977a );
 a46984a <=( (not A203)  and  (not A202) );
 a46987a <=( (not A235)  and  (not A234) );
 a46988a <=( a46987a  and  a46984a );
 a46989a <=( a46988a  and  a46981a );
 a46992a <=( A265  and  (not A236) );
 a46995a <=( (not A267)  and  A266 );
 a46996a <=( a46995a  and  a46992a );
 a46999a <=( (not A300)  and  (not A268) );
 a47002a <=( (not A302)  and  (not A301) );
 a47003a <=( a47002a  and  a46999a );
 a47004a <=( a47003a  and  a46996a );
 a47007a <=( (not A167)  and  A170 );
 a47010a <=( (not A201)  and  A166 );
 a47011a <=( a47010a  and  a47007a );
 a47014a <=( (not A203)  and  (not A202) );
 a47017a <=( (not A235)  and  (not A234) );
 a47018a <=( a47017a  and  a47014a );
 a47019a <=( a47018a  and  a47011a );
 a47022a <=( A265  and  (not A236) );
 a47025a <=( (not A267)  and  A266 );
 a47026a <=( a47025a  and  a47022a );
 a47029a <=( (not A298)  and  (not A268) );
 a47032a <=( (not A301)  and  (not A299) );
 a47033a <=( a47032a  and  a47029a );
 a47034a <=( a47033a  and  a47026a );
 a47037a <=( (not A167)  and  A170 );
 a47040a <=( (not A201)  and  A166 );
 a47041a <=( a47040a  and  a47037a );
 a47044a <=( (not A203)  and  (not A202) );
 a47047a <=( (not A235)  and  (not A234) );
 a47048a <=( a47047a  and  a47044a );
 a47049a <=( a47048a  and  a47041a );
 a47052a <=( (not A265)  and  (not A236) );
 a47055a <=( (not A268)  and  (not A266) );
 a47056a <=( a47055a  and  a47052a );
 a47059a <=( A299  and  A298 );
 a47062a <=( (not A301)  and  (not A300) );
 a47063a <=( a47062a  and  a47059a );
 a47064a <=( a47063a  and  a47056a );
 a47067a <=( (not A167)  and  A170 );
 a47070a <=( (not A201)  and  A166 );
 a47071a <=( a47070a  and  a47067a );
 a47074a <=( (not A203)  and  (not A202) );
 a47077a <=( A233  and  A232 );
 a47078a <=( a47077a  and  a47074a );
 a47079a <=( a47078a  and  a47071a );
 a47082a <=( (not A235)  and  (not A234) );
 a47085a <=( (not A268)  and  (not A267) );
 a47086a <=( a47085a  and  a47082a );
 a47089a <=( (not A300)  and  (not A269) );
 a47092a <=( (not A302)  and  (not A301) );
 a47093a <=( a47092a  and  a47089a );
 a47094a <=( a47093a  and  a47086a );
 a47097a <=( (not A167)  and  A170 );
 a47100a <=( (not A201)  and  A166 );
 a47101a <=( a47100a  and  a47097a );
 a47104a <=( (not A203)  and  (not A202) );
 a47107a <=( A233  and  A232 );
 a47108a <=( a47107a  and  a47104a );
 a47109a <=( a47108a  and  a47101a );
 a47112a <=( (not A235)  and  (not A234) );
 a47115a <=( (not A268)  and  (not A267) );
 a47116a <=( a47115a  and  a47112a );
 a47119a <=( (not A298)  and  (not A269) );
 a47122a <=( (not A301)  and  (not A299) );
 a47123a <=( a47122a  and  a47119a );
 a47124a <=( a47123a  and  a47116a );
 a47127a <=( (not A167)  and  A170 );
 a47130a <=( (not A201)  and  A166 );
 a47131a <=( a47130a  and  a47127a );
 a47134a <=( (not A203)  and  (not A202) );
 a47137a <=( A233  and  A232 );
 a47138a <=( a47137a  and  a47134a );
 a47139a <=( a47138a  and  a47131a );
 a47142a <=( (not A235)  and  (not A234) );
 a47145a <=( (not A266)  and  (not A265) );
 a47146a <=( a47145a  and  a47142a );
 a47149a <=( (not A300)  and  (not A268) );
 a47152a <=( (not A302)  and  (not A301) );
 a47153a <=( a47152a  and  a47149a );
 a47154a <=( a47153a  and  a47146a );
 a47157a <=( (not A167)  and  A170 );
 a47160a <=( (not A201)  and  A166 );
 a47161a <=( a47160a  and  a47157a );
 a47164a <=( (not A203)  and  (not A202) );
 a47167a <=( A233  and  A232 );
 a47168a <=( a47167a  and  a47164a );
 a47169a <=( a47168a  and  a47161a );
 a47172a <=( (not A235)  and  (not A234) );
 a47175a <=( (not A266)  and  (not A265) );
 a47176a <=( a47175a  and  a47172a );
 a47179a <=( (not A298)  and  (not A268) );
 a47182a <=( (not A301)  and  (not A299) );
 a47183a <=( a47182a  and  a47179a );
 a47184a <=( a47183a  and  a47176a );
 a47187a <=( (not A167)  and  A170 );
 a47190a <=( (not A201)  and  A166 );
 a47191a <=( a47190a  and  a47187a );
 a47194a <=( (not A203)  and  (not A202) );
 a47197a <=( (not A233)  and  (not A232) );
 a47198a <=( a47197a  and  a47194a );
 a47199a <=( a47198a  and  a47191a );
 a47202a <=( (not A267)  and  (not A235) );
 a47205a <=( (not A269)  and  (not A268) );
 a47206a <=( a47205a  and  a47202a );
 a47209a <=( A299  and  A298 );
 a47212a <=( (not A301)  and  (not A300) );
 a47213a <=( a47212a  and  a47209a );
 a47214a <=( a47213a  and  a47206a );
 a47217a <=( (not A167)  and  A170 );
 a47220a <=( (not A201)  and  A166 );
 a47221a <=( a47220a  and  a47217a );
 a47224a <=( (not A203)  and  (not A202) );
 a47227a <=( (not A233)  and  (not A232) );
 a47228a <=( a47227a  and  a47224a );
 a47229a <=( a47228a  and  a47221a );
 a47232a <=( A265  and  (not A235) );
 a47235a <=( (not A267)  and  A266 );
 a47236a <=( a47235a  and  a47232a );
 a47239a <=( (not A300)  and  (not A268) );
 a47242a <=( (not A302)  and  (not A301) );
 a47243a <=( a47242a  and  a47239a );
 a47244a <=( a47243a  and  a47236a );
 a47247a <=( (not A167)  and  A170 );
 a47250a <=( (not A201)  and  A166 );
 a47251a <=( a47250a  and  a47247a );
 a47254a <=( (not A203)  and  (not A202) );
 a47257a <=( (not A233)  and  (not A232) );
 a47258a <=( a47257a  and  a47254a );
 a47259a <=( a47258a  and  a47251a );
 a47262a <=( A265  and  (not A235) );
 a47265a <=( (not A267)  and  A266 );
 a47266a <=( a47265a  and  a47262a );
 a47269a <=( (not A298)  and  (not A268) );
 a47272a <=( (not A301)  and  (not A299) );
 a47273a <=( a47272a  and  a47269a );
 a47274a <=( a47273a  and  a47266a );
 a47277a <=( (not A167)  and  A170 );
 a47280a <=( (not A201)  and  A166 );
 a47281a <=( a47280a  and  a47277a );
 a47284a <=( (not A203)  and  (not A202) );
 a47287a <=( (not A233)  and  (not A232) );
 a47288a <=( a47287a  and  a47284a );
 a47289a <=( a47288a  and  a47281a );
 a47292a <=( (not A265)  and  (not A235) );
 a47295a <=( (not A268)  and  (not A266) );
 a47296a <=( a47295a  and  a47292a );
 a47299a <=( A299  and  A298 );
 a47302a <=( (not A301)  and  (not A300) );
 a47303a <=( a47302a  and  a47299a );
 a47304a <=( a47303a  and  a47296a );
 a47307a <=( (not A167)  and  A170 );
 a47310a <=( A199  and  A166 );
 a47311a <=( a47310a  and  a47307a );
 a47314a <=( (not A201)  and  A200 );
 a47317a <=( (not A234)  and  (not A202) );
 a47318a <=( a47317a  and  a47314a );
 a47319a <=( a47318a  and  a47311a );
 a47322a <=( (not A236)  and  (not A235) );
 a47325a <=( (not A268)  and  (not A267) );
 a47326a <=( a47325a  and  a47322a );
 a47329a <=( (not A300)  and  (not A269) );
 a47332a <=( (not A302)  and  (not A301) );
 a47333a <=( a47332a  and  a47329a );
 a47334a <=( a47333a  and  a47326a );
 a47337a <=( (not A167)  and  A170 );
 a47340a <=( A199  and  A166 );
 a47341a <=( a47340a  and  a47337a );
 a47344a <=( (not A201)  and  A200 );
 a47347a <=( (not A234)  and  (not A202) );
 a47348a <=( a47347a  and  a47344a );
 a47349a <=( a47348a  and  a47341a );
 a47352a <=( (not A236)  and  (not A235) );
 a47355a <=( (not A268)  and  (not A267) );
 a47356a <=( a47355a  and  a47352a );
 a47359a <=( (not A298)  and  (not A269) );
 a47362a <=( (not A301)  and  (not A299) );
 a47363a <=( a47362a  and  a47359a );
 a47364a <=( a47363a  and  a47356a );
 a47367a <=( (not A167)  and  A170 );
 a47370a <=( A199  and  A166 );
 a47371a <=( a47370a  and  a47367a );
 a47374a <=( (not A201)  and  A200 );
 a47377a <=( (not A234)  and  (not A202) );
 a47378a <=( a47377a  and  a47374a );
 a47379a <=( a47378a  and  a47371a );
 a47382a <=( (not A236)  and  (not A235) );
 a47385a <=( (not A266)  and  (not A265) );
 a47386a <=( a47385a  and  a47382a );
 a47389a <=( (not A300)  and  (not A268) );
 a47392a <=( (not A302)  and  (not A301) );
 a47393a <=( a47392a  and  a47389a );
 a47394a <=( a47393a  and  a47386a );
 a47397a <=( (not A167)  and  A170 );
 a47400a <=( A199  and  A166 );
 a47401a <=( a47400a  and  a47397a );
 a47404a <=( (not A201)  and  A200 );
 a47407a <=( (not A234)  and  (not A202) );
 a47408a <=( a47407a  and  a47404a );
 a47409a <=( a47408a  and  a47401a );
 a47412a <=( (not A236)  and  (not A235) );
 a47415a <=( (not A266)  and  (not A265) );
 a47416a <=( a47415a  and  a47412a );
 a47419a <=( (not A298)  and  (not A268) );
 a47422a <=( (not A301)  and  (not A299) );
 a47423a <=( a47422a  and  a47419a );
 a47424a <=( a47423a  and  a47416a );
 a47427a <=( (not A167)  and  A170 );
 a47430a <=( A199  and  A166 );
 a47431a <=( a47430a  and  a47427a );
 a47434a <=( (not A201)  and  A200 );
 a47437a <=( (not A232)  and  (not A202) );
 a47438a <=( a47437a  and  a47434a );
 a47439a <=( a47438a  and  a47431a );
 a47442a <=( (not A235)  and  (not A233) );
 a47445a <=( (not A268)  and  (not A267) );
 a47446a <=( a47445a  and  a47442a );
 a47449a <=( (not A300)  and  (not A269) );
 a47452a <=( (not A302)  and  (not A301) );
 a47453a <=( a47452a  and  a47449a );
 a47454a <=( a47453a  and  a47446a );
 a47457a <=( (not A167)  and  A170 );
 a47460a <=( A199  and  A166 );
 a47461a <=( a47460a  and  a47457a );
 a47464a <=( (not A201)  and  A200 );
 a47467a <=( (not A232)  and  (not A202) );
 a47468a <=( a47467a  and  a47464a );
 a47469a <=( a47468a  and  a47461a );
 a47472a <=( (not A235)  and  (not A233) );
 a47475a <=( (not A268)  and  (not A267) );
 a47476a <=( a47475a  and  a47472a );
 a47479a <=( (not A298)  and  (not A269) );
 a47482a <=( (not A301)  and  (not A299) );
 a47483a <=( a47482a  and  a47479a );
 a47484a <=( a47483a  and  a47476a );
 a47487a <=( (not A167)  and  A170 );
 a47490a <=( A199  and  A166 );
 a47491a <=( a47490a  and  a47487a );
 a47494a <=( (not A201)  and  A200 );
 a47497a <=( (not A232)  and  (not A202) );
 a47498a <=( a47497a  and  a47494a );
 a47499a <=( a47498a  and  a47491a );
 a47502a <=( (not A235)  and  (not A233) );
 a47505a <=( (not A266)  and  (not A265) );
 a47506a <=( a47505a  and  a47502a );
 a47509a <=( (not A300)  and  (not A268) );
 a47512a <=( (not A302)  and  (not A301) );
 a47513a <=( a47512a  and  a47509a );
 a47514a <=( a47513a  and  a47506a );
 a47517a <=( (not A167)  and  A170 );
 a47520a <=( A199  and  A166 );
 a47521a <=( a47520a  and  a47517a );
 a47524a <=( (not A201)  and  A200 );
 a47527a <=( (not A232)  and  (not A202) );
 a47528a <=( a47527a  and  a47524a );
 a47529a <=( a47528a  and  a47521a );
 a47532a <=( (not A235)  and  (not A233) );
 a47535a <=( (not A266)  and  (not A265) );
 a47536a <=( a47535a  and  a47532a );
 a47539a <=( (not A298)  and  (not A268) );
 a47542a <=( (not A301)  and  (not A299) );
 a47543a <=( a47542a  and  a47539a );
 a47544a <=( a47543a  and  a47536a );
 a47547a <=( (not A167)  and  A170 );
 a47550a <=( (not A199)  and  A166 );
 a47551a <=( a47550a  and  a47547a );
 a47554a <=( (not A202)  and  (not A200) );
 a47557a <=( (not A235)  and  (not A234) );
 a47558a <=( a47557a  and  a47554a );
 a47559a <=( a47558a  and  a47551a );
 a47562a <=( (not A267)  and  (not A236) );
 a47565a <=( (not A269)  and  (not A268) );
 a47566a <=( a47565a  and  a47562a );
 a47569a <=( A299  and  A298 );
 a47572a <=( (not A301)  and  (not A300) );
 a47573a <=( a47572a  and  a47569a );
 a47574a <=( a47573a  and  a47566a );
 a47577a <=( (not A167)  and  A170 );
 a47580a <=( (not A199)  and  A166 );
 a47581a <=( a47580a  and  a47577a );
 a47584a <=( (not A202)  and  (not A200) );
 a47587a <=( (not A235)  and  (not A234) );
 a47588a <=( a47587a  and  a47584a );
 a47589a <=( a47588a  and  a47581a );
 a47592a <=( A265  and  (not A236) );
 a47595a <=( (not A267)  and  A266 );
 a47596a <=( a47595a  and  a47592a );
 a47599a <=( (not A300)  and  (not A268) );
 a47602a <=( (not A302)  and  (not A301) );
 a47603a <=( a47602a  and  a47599a );
 a47604a <=( a47603a  and  a47596a );
 a47607a <=( (not A167)  and  A170 );
 a47610a <=( (not A199)  and  A166 );
 a47611a <=( a47610a  and  a47607a );
 a47614a <=( (not A202)  and  (not A200) );
 a47617a <=( (not A235)  and  (not A234) );
 a47618a <=( a47617a  and  a47614a );
 a47619a <=( a47618a  and  a47611a );
 a47622a <=( A265  and  (not A236) );
 a47625a <=( (not A267)  and  A266 );
 a47626a <=( a47625a  and  a47622a );
 a47629a <=( (not A298)  and  (not A268) );
 a47632a <=( (not A301)  and  (not A299) );
 a47633a <=( a47632a  and  a47629a );
 a47634a <=( a47633a  and  a47626a );
 a47637a <=( (not A167)  and  A170 );
 a47640a <=( (not A199)  and  A166 );
 a47641a <=( a47640a  and  a47637a );
 a47644a <=( (not A202)  and  (not A200) );
 a47647a <=( (not A235)  and  (not A234) );
 a47648a <=( a47647a  and  a47644a );
 a47649a <=( a47648a  and  a47641a );
 a47652a <=( (not A265)  and  (not A236) );
 a47655a <=( (not A268)  and  (not A266) );
 a47656a <=( a47655a  and  a47652a );
 a47659a <=( A299  and  A298 );
 a47662a <=( (not A301)  and  (not A300) );
 a47663a <=( a47662a  and  a47659a );
 a47664a <=( a47663a  and  a47656a );
 a47667a <=( (not A167)  and  A170 );
 a47670a <=( (not A199)  and  A166 );
 a47671a <=( a47670a  and  a47667a );
 a47674a <=( (not A202)  and  (not A200) );
 a47677a <=( A233  and  A232 );
 a47678a <=( a47677a  and  a47674a );
 a47679a <=( a47678a  and  a47671a );
 a47682a <=( (not A235)  and  (not A234) );
 a47685a <=( (not A268)  and  (not A267) );
 a47686a <=( a47685a  and  a47682a );
 a47689a <=( (not A300)  and  (not A269) );
 a47692a <=( (not A302)  and  (not A301) );
 a47693a <=( a47692a  and  a47689a );
 a47694a <=( a47693a  and  a47686a );
 a47697a <=( (not A167)  and  A170 );
 a47700a <=( (not A199)  and  A166 );
 a47701a <=( a47700a  and  a47697a );
 a47704a <=( (not A202)  and  (not A200) );
 a47707a <=( A233  and  A232 );
 a47708a <=( a47707a  and  a47704a );
 a47709a <=( a47708a  and  a47701a );
 a47712a <=( (not A235)  and  (not A234) );
 a47715a <=( (not A268)  and  (not A267) );
 a47716a <=( a47715a  and  a47712a );
 a47719a <=( (not A298)  and  (not A269) );
 a47722a <=( (not A301)  and  (not A299) );
 a47723a <=( a47722a  and  a47719a );
 a47724a <=( a47723a  and  a47716a );
 a47727a <=( (not A167)  and  A170 );
 a47730a <=( (not A199)  and  A166 );
 a47731a <=( a47730a  and  a47727a );
 a47734a <=( (not A202)  and  (not A200) );
 a47737a <=( A233  and  A232 );
 a47738a <=( a47737a  and  a47734a );
 a47739a <=( a47738a  and  a47731a );
 a47742a <=( (not A235)  and  (not A234) );
 a47745a <=( (not A266)  and  (not A265) );
 a47746a <=( a47745a  and  a47742a );
 a47749a <=( (not A300)  and  (not A268) );
 a47752a <=( (not A302)  and  (not A301) );
 a47753a <=( a47752a  and  a47749a );
 a47754a <=( a47753a  and  a47746a );
 a47757a <=( (not A167)  and  A170 );
 a47760a <=( (not A199)  and  A166 );
 a47761a <=( a47760a  and  a47757a );
 a47764a <=( (not A202)  and  (not A200) );
 a47767a <=( A233  and  A232 );
 a47768a <=( a47767a  and  a47764a );
 a47769a <=( a47768a  and  a47761a );
 a47772a <=( (not A235)  and  (not A234) );
 a47775a <=( (not A266)  and  (not A265) );
 a47776a <=( a47775a  and  a47772a );
 a47779a <=( (not A298)  and  (not A268) );
 a47782a <=( (not A301)  and  (not A299) );
 a47783a <=( a47782a  and  a47779a );
 a47784a <=( a47783a  and  a47776a );
 a47787a <=( (not A167)  and  A170 );
 a47790a <=( (not A199)  and  A166 );
 a47791a <=( a47790a  and  a47787a );
 a47794a <=( (not A202)  and  (not A200) );
 a47797a <=( (not A233)  and  (not A232) );
 a47798a <=( a47797a  and  a47794a );
 a47799a <=( a47798a  and  a47791a );
 a47802a <=( (not A267)  and  (not A235) );
 a47805a <=( (not A269)  and  (not A268) );
 a47806a <=( a47805a  and  a47802a );
 a47809a <=( A299  and  A298 );
 a47812a <=( (not A301)  and  (not A300) );
 a47813a <=( a47812a  and  a47809a );
 a47814a <=( a47813a  and  a47806a );
 a47817a <=( (not A167)  and  A170 );
 a47820a <=( (not A199)  and  A166 );
 a47821a <=( a47820a  and  a47817a );
 a47824a <=( (not A202)  and  (not A200) );
 a47827a <=( (not A233)  and  (not A232) );
 a47828a <=( a47827a  and  a47824a );
 a47829a <=( a47828a  and  a47821a );
 a47832a <=( A265  and  (not A235) );
 a47835a <=( (not A267)  and  A266 );
 a47836a <=( a47835a  and  a47832a );
 a47839a <=( (not A300)  and  (not A268) );
 a47842a <=( (not A302)  and  (not A301) );
 a47843a <=( a47842a  and  a47839a );
 a47844a <=( a47843a  and  a47836a );
 a47847a <=( (not A167)  and  A170 );
 a47850a <=( (not A199)  and  A166 );
 a47851a <=( a47850a  and  a47847a );
 a47854a <=( (not A202)  and  (not A200) );
 a47857a <=( (not A233)  and  (not A232) );
 a47858a <=( a47857a  and  a47854a );
 a47859a <=( a47858a  and  a47851a );
 a47862a <=( A265  and  (not A235) );
 a47865a <=( (not A267)  and  A266 );
 a47866a <=( a47865a  and  a47862a );
 a47869a <=( (not A298)  and  (not A268) );
 a47872a <=( (not A301)  and  (not A299) );
 a47873a <=( a47872a  and  a47869a );
 a47874a <=( a47873a  and  a47866a );
 a47877a <=( (not A167)  and  A170 );
 a47880a <=( (not A199)  and  A166 );
 a47881a <=( a47880a  and  a47877a );
 a47884a <=( (not A202)  and  (not A200) );
 a47887a <=( (not A233)  and  (not A232) );
 a47888a <=( a47887a  and  a47884a );
 a47889a <=( a47888a  and  a47881a );
 a47892a <=( (not A265)  and  (not A235) );
 a47895a <=( (not A268)  and  (not A266) );
 a47896a <=( a47895a  and  a47892a );
 a47899a <=( A299  and  A298 );
 a47902a <=( (not A301)  and  (not A300) );
 a47903a <=( a47902a  and  a47899a );
 a47904a <=( a47903a  and  a47896a );
 a47907a <=( (not A201)  and  A169 );
 a47910a <=( (not A203)  and  (not A202) );
 a47911a <=( a47910a  and  a47907a );
 a47914a <=( A233  and  A232 );
 a47917a <=( (not A235)  and  (not A234) );
 a47918a <=( a47917a  and  a47914a );
 a47919a <=( a47918a  and  a47911a );
 a47922a <=( A266  and  A265 );
 a47925a <=( (not A268)  and  (not A267) );
 a47926a <=( a47925a  and  a47922a );
 a47929a <=( A299  and  A298 );
 a47932a <=( (not A301)  and  (not A300) );
 a47933a <=( a47932a  and  a47929a );
 a47934a <=( a47933a  and  a47926a );
 a47937a <=( A199  and  A169 );
 a47940a <=( (not A201)  and  A200 );
 a47941a <=( a47940a  and  a47937a );
 a47944a <=( (not A234)  and  (not A202) );
 a47947a <=( (not A236)  and  (not A235) );
 a47948a <=( a47947a  and  a47944a );
 a47949a <=( a47948a  and  a47941a );
 a47952a <=( A266  and  A265 );
 a47955a <=( (not A268)  and  (not A267) );
 a47956a <=( a47955a  and  a47952a );
 a47959a <=( A299  and  A298 );
 a47962a <=( (not A301)  and  (not A300) );
 a47963a <=( a47962a  and  a47959a );
 a47964a <=( a47963a  and  a47956a );
 a47967a <=( A199  and  A169 );
 a47970a <=( (not A201)  and  A200 );
 a47971a <=( a47970a  and  a47967a );
 a47974a <=( A232  and  (not A202) );
 a47977a <=( (not A234)  and  A233 );
 a47978a <=( a47977a  and  a47974a );
 a47979a <=( a47978a  and  a47971a );
 a47982a <=( (not A267)  and  (not A235) );
 a47985a <=( (not A269)  and  (not A268) );
 a47986a <=( a47985a  and  a47982a );
 a47989a <=( A299  and  A298 );
 a47992a <=( (not A301)  and  (not A300) );
 a47993a <=( a47992a  and  a47989a );
 a47994a <=( a47993a  and  a47986a );
 a47997a <=( A199  and  A169 );
 a48000a <=( (not A201)  and  A200 );
 a48001a <=( a48000a  and  a47997a );
 a48004a <=( A232  and  (not A202) );
 a48007a <=( (not A234)  and  A233 );
 a48008a <=( a48007a  and  a48004a );
 a48009a <=( a48008a  and  a48001a );
 a48012a <=( A265  and  (not A235) );
 a48015a <=( (not A267)  and  A266 );
 a48016a <=( a48015a  and  a48012a );
 a48019a <=( (not A300)  and  (not A268) );
 a48022a <=( (not A302)  and  (not A301) );
 a48023a <=( a48022a  and  a48019a );
 a48024a <=( a48023a  and  a48016a );
 a48027a <=( A199  and  A169 );
 a48030a <=( (not A201)  and  A200 );
 a48031a <=( a48030a  and  a48027a );
 a48034a <=( A232  and  (not A202) );
 a48037a <=( (not A234)  and  A233 );
 a48038a <=( a48037a  and  a48034a );
 a48039a <=( a48038a  and  a48031a );
 a48042a <=( A265  and  (not A235) );
 a48045a <=( (not A267)  and  A266 );
 a48046a <=( a48045a  and  a48042a );
 a48049a <=( (not A298)  and  (not A268) );
 a48052a <=( (not A301)  and  (not A299) );
 a48053a <=( a48052a  and  a48049a );
 a48054a <=( a48053a  and  a48046a );
 a48057a <=( A199  and  A169 );
 a48060a <=( (not A201)  and  A200 );
 a48061a <=( a48060a  and  a48057a );
 a48064a <=( A232  and  (not A202) );
 a48067a <=( (not A234)  and  A233 );
 a48068a <=( a48067a  and  a48064a );
 a48069a <=( a48068a  and  a48061a );
 a48072a <=( (not A265)  and  (not A235) );
 a48075a <=( (not A268)  and  (not A266) );
 a48076a <=( a48075a  and  a48072a );
 a48079a <=( A299  and  A298 );
 a48082a <=( (not A301)  and  (not A300) );
 a48083a <=( a48082a  and  a48079a );
 a48084a <=( a48083a  and  a48076a );
 a48087a <=( A199  and  A169 );
 a48090a <=( (not A201)  and  A200 );
 a48091a <=( a48090a  and  a48087a );
 a48094a <=( (not A232)  and  (not A202) );
 a48097a <=( (not A235)  and  (not A233) );
 a48098a <=( a48097a  and  a48094a );
 a48099a <=( a48098a  and  a48091a );
 a48102a <=( A266  and  A265 );
 a48105a <=( (not A268)  and  (not A267) );
 a48106a <=( a48105a  and  a48102a );
 a48109a <=( A299  and  A298 );
 a48112a <=( (not A301)  and  (not A300) );
 a48113a <=( a48112a  and  a48109a );
 a48114a <=( a48113a  and  a48106a );
 a48117a <=( (not A199)  and  A169 );
 a48120a <=( (not A202)  and  (not A200) );
 a48121a <=( a48120a  and  a48117a );
 a48124a <=( A233  and  A232 );
 a48127a <=( (not A235)  and  (not A234) );
 a48128a <=( a48127a  and  a48124a );
 a48129a <=( a48128a  and  a48121a );
 a48132a <=( A266  and  A265 );
 a48135a <=( (not A268)  and  (not A267) );
 a48136a <=( a48135a  and  a48132a );
 a48139a <=( A299  and  A298 );
 a48142a <=( (not A301)  and  (not A300) );
 a48143a <=( a48142a  and  a48139a );
 a48144a <=( a48143a  and  a48136a );
 a48147a <=( (not A167)  and  (not A169) );
 a48150a <=( A202  and  (not A166) );
 a48151a <=( a48150a  and  a48147a );
 a48154a <=( A233  and  A232 );
 a48157a <=( (not A235)  and  (not A234) );
 a48158a <=( a48157a  and  a48154a );
 a48159a <=( a48158a  and  a48151a );
 a48162a <=( A266  and  A265 );
 a48165a <=( (not A268)  and  (not A267) );
 a48166a <=( a48165a  and  a48162a );
 a48169a <=( A299  and  A298 );
 a48172a <=( (not A301)  and  (not A300) );
 a48173a <=( a48172a  and  a48169a );
 a48174a <=( a48173a  and  a48166a );
 a48177a <=( (not A167)  and  (not A169) );
 a48180a <=( A199  and  (not A166) );
 a48181a <=( a48180a  and  a48177a );
 a48184a <=( (not A234)  and  A201 );
 a48187a <=( (not A236)  and  (not A235) );
 a48188a <=( a48187a  and  a48184a );
 a48189a <=( a48188a  and  a48181a );
 a48192a <=( A266  and  A265 );
 a48195a <=( (not A268)  and  (not A267) );
 a48196a <=( a48195a  and  a48192a );
 a48199a <=( A299  and  A298 );
 a48202a <=( (not A301)  and  (not A300) );
 a48203a <=( a48202a  and  a48199a );
 a48204a <=( a48203a  and  a48196a );
 a48207a <=( (not A167)  and  (not A169) );
 a48210a <=( A199  and  (not A166) );
 a48211a <=( a48210a  and  a48207a );
 a48214a <=( A232  and  A201 );
 a48217a <=( (not A234)  and  A233 );
 a48218a <=( a48217a  and  a48214a );
 a48219a <=( a48218a  and  a48211a );
 a48222a <=( (not A267)  and  (not A235) );
 a48225a <=( (not A269)  and  (not A268) );
 a48226a <=( a48225a  and  a48222a );
 a48229a <=( A299  and  A298 );
 a48232a <=( (not A301)  and  (not A300) );
 a48233a <=( a48232a  and  a48229a );
 a48234a <=( a48233a  and  a48226a );
 a48237a <=( (not A167)  and  (not A169) );
 a48240a <=( A199  and  (not A166) );
 a48241a <=( a48240a  and  a48237a );
 a48244a <=( A232  and  A201 );
 a48247a <=( (not A234)  and  A233 );
 a48248a <=( a48247a  and  a48244a );
 a48249a <=( a48248a  and  a48241a );
 a48252a <=( A265  and  (not A235) );
 a48255a <=( (not A267)  and  A266 );
 a48256a <=( a48255a  and  a48252a );
 a48259a <=( (not A300)  and  (not A268) );
 a48262a <=( (not A302)  and  (not A301) );
 a48263a <=( a48262a  and  a48259a );
 a48264a <=( a48263a  and  a48256a );
 a48267a <=( (not A167)  and  (not A169) );
 a48270a <=( A199  and  (not A166) );
 a48271a <=( a48270a  and  a48267a );
 a48274a <=( A232  and  A201 );
 a48277a <=( (not A234)  and  A233 );
 a48278a <=( a48277a  and  a48274a );
 a48279a <=( a48278a  and  a48271a );
 a48282a <=( A265  and  (not A235) );
 a48285a <=( (not A267)  and  A266 );
 a48286a <=( a48285a  and  a48282a );
 a48289a <=( (not A298)  and  (not A268) );
 a48292a <=( (not A301)  and  (not A299) );
 a48293a <=( a48292a  and  a48289a );
 a48294a <=( a48293a  and  a48286a );
 a48297a <=( (not A167)  and  (not A169) );
 a48300a <=( A199  and  (not A166) );
 a48301a <=( a48300a  and  a48297a );
 a48304a <=( A232  and  A201 );
 a48307a <=( (not A234)  and  A233 );
 a48308a <=( a48307a  and  a48304a );
 a48309a <=( a48308a  and  a48301a );
 a48312a <=( (not A265)  and  (not A235) );
 a48315a <=( (not A268)  and  (not A266) );
 a48316a <=( a48315a  and  a48312a );
 a48319a <=( A299  and  A298 );
 a48322a <=( (not A301)  and  (not A300) );
 a48323a <=( a48322a  and  a48319a );
 a48324a <=( a48323a  and  a48316a );
 a48327a <=( (not A167)  and  (not A169) );
 a48330a <=( A199  and  (not A166) );
 a48331a <=( a48330a  and  a48327a );
 a48334a <=( (not A232)  and  A201 );
 a48337a <=( (not A235)  and  (not A233) );
 a48338a <=( a48337a  and  a48334a );
 a48339a <=( a48338a  and  a48331a );
 a48342a <=( A266  and  A265 );
 a48345a <=( (not A268)  and  (not A267) );
 a48346a <=( a48345a  and  a48342a );
 a48349a <=( A299  and  A298 );
 a48352a <=( (not A301)  and  (not A300) );
 a48353a <=( a48352a  and  a48349a );
 a48354a <=( a48353a  and  a48346a );
 a48357a <=( (not A167)  and  (not A169) );
 a48360a <=( A200  and  (not A166) );
 a48361a <=( a48360a  and  a48357a );
 a48364a <=( (not A234)  and  A201 );
 a48367a <=( (not A236)  and  (not A235) );
 a48368a <=( a48367a  and  a48364a );
 a48369a <=( a48368a  and  a48361a );
 a48372a <=( A266  and  A265 );
 a48375a <=( (not A268)  and  (not A267) );
 a48376a <=( a48375a  and  a48372a );
 a48379a <=( A299  and  A298 );
 a48382a <=( (not A301)  and  (not A300) );
 a48383a <=( a48382a  and  a48379a );
 a48384a <=( a48383a  and  a48376a );
 a48387a <=( (not A167)  and  (not A169) );
 a48390a <=( A200  and  (not A166) );
 a48391a <=( a48390a  and  a48387a );
 a48394a <=( A232  and  A201 );
 a48397a <=( (not A234)  and  A233 );
 a48398a <=( a48397a  and  a48394a );
 a48399a <=( a48398a  and  a48391a );
 a48402a <=( (not A267)  and  (not A235) );
 a48405a <=( (not A269)  and  (not A268) );
 a48406a <=( a48405a  and  a48402a );
 a48409a <=( A299  and  A298 );
 a48412a <=( (not A301)  and  (not A300) );
 a48413a <=( a48412a  and  a48409a );
 a48414a <=( a48413a  and  a48406a );
 a48417a <=( (not A167)  and  (not A169) );
 a48420a <=( A200  and  (not A166) );
 a48421a <=( a48420a  and  a48417a );
 a48424a <=( A232  and  A201 );
 a48427a <=( (not A234)  and  A233 );
 a48428a <=( a48427a  and  a48424a );
 a48429a <=( a48428a  and  a48421a );
 a48432a <=( A265  and  (not A235) );
 a48435a <=( (not A267)  and  A266 );
 a48436a <=( a48435a  and  a48432a );
 a48439a <=( (not A300)  and  (not A268) );
 a48442a <=( (not A302)  and  (not A301) );
 a48443a <=( a48442a  and  a48439a );
 a48444a <=( a48443a  and  a48436a );
 a48447a <=( (not A167)  and  (not A169) );
 a48450a <=( A200  and  (not A166) );
 a48451a <=( a48450a  and  a48447a );
 a48454a <=( A232  and  A201 );
 a48457a <=( (not A234)  and  A233 );
 a48458a <=( a48457a  and  a48454a );
 a48459a <=( a48458a  and  a48451a );
 a48462a <=( A265  and  (not A235) );
 a48465a <=( (not A267)  and  A266 );
 a48466a <=( a48465a  and  a48462a );
 a48469a <=( (not A298)  and  (not A268) );
 a48472a <=( (not A301)  and  (not A299) );
 a48473a <=( a48472a  and  a48469a );
 a48474a <=( a48473a  and  a48466a );
 a48477a <=( (not A167)  and  (not A169) );
 a48480a <=( A200  and  (not A166) );
 a48481a <=( a48480a  and  a48477a );
 a48484a <=( A232  and  A201 );
 a48487a <=( (not A234)  and  A233 );
 a48488a <=( a48487a  and  a48484a );
 a48489a <=( a48488a  and  a48481a );
 a48492a <=( (not A265)  and  (not A235) );
 a48495a <=( (not A268)  and  (not A266) );
 a48496a <=( a48495a  and  a48492a );
 a48499a <=( A299  and  A298 );
 a48502a <=( (not A301)  and  (not A300) );
 a48503a <=( a48502a  and  a48499a );
 a48504a <=( a48503a  and  a48496a );
 a48507a <=( (not A167)  and  (not A169) );
 a48510a <=( A200  and  (not A166) );
 a48511a <=( a48510a  and  a48507a );
 a48514a <=( (not A232)  and  A201 );
 a48517a <=( (not A235)  and  (not A233) );
 a48518a <=( a48517a  and  a48514a );
 a48519a <=( a48518a  and  a48511a );
 a48522a <=( A266  and  A265 );
 a48525a <=( (not A268)  and  (not A267) );
 a48526a <=( a48525a  and  a48522a );
 a48529a <=( A299  and  A298 );
 a48532a <=( (not A301)  and  (not A300) );
 a48533a <=( a48532a  and  a48529a );
 a48534a <=( a48533a  and  a48526a );
 a48537a <=( (not A167)  and  (not A169) );
 a48540a <=( (not A199)  and  (not A166) );
 a48541a <=( a48540a  and  a48537a );
 a48544a <=( A203  and  A200 );
 a48547a <=( (not A235)  and  (not A234) );
 a48548a <=( a48547a  and  a48544a );
 a48549a <=( a48548a  and  a48541a );
 a48552a <=( (not A267)  and  (not A236) );
 a48555a <=( (not A269)  and  (not A268) );
 a48556a <=( a48555a  and  a48552a );
 a48559a <=( A299  and  A298 );
 a48562a <=( (not A301)  and  (not A300) );
 a48563a <=( a48562a  and  a48559a );
 a48564a <=( a48563a  and  a48556a );
 a48567a <=( (not A167)  and  (not A169) );
 a48570a <=( (not A199)  and  (not A166) );
 a48571a <=( a48570a  and  a48567a );
 a48574a <=( A203  and  A200 );
 a48577a <=( (not A235)  and  (not A234) );
 a48578a <=( a48577a  and  a48574a );
 a48579a <=( a48578a  and  a48571a );
 a48582a <=( A265  and  (not A236) );
 a48585a <=( (not A267)  and  A266 );
 a48586a <=( a48585a  and  a48582a );
 a48589a <=( (not A300)  and  (not A268) );
 a48592a <=( (not A302)  and  (not A301) );
 a48593a <=( a48592a  and  a48589a );
 a48594a <=( a48593a  and  a48586a );
 a48597a <=( (not A167)  and  (not A169) );
 a48600a <=( (not A199)  and  (not A166) );
 a48601a <=( a48600a  and  a48597a );
 a48604a <=( A203  and  A200 );
 a48607a <=( (not A235)  and  (not A234) );
 a48608a <=( a48607a  and  a48604a );
 a48609a <=( a48608a  and  a48601a );
 a48612a <=( A265  and  (not A236) );
 a48615a <=( (not A267)  and  A266 );
 a48616a <=( a48615a  and  a48612a );
 a48619a <=( (not A298)  and  (not A268) );
 a48622a <=( (not A301)  and  (not A299) );
 a48623a <=( a48622a  and  a48619a );
 a48624a <=( a48623a  and  a48616a );
 a48627a <=( (not A167)  and  (not A169) );
 a48630a <=( (not A199)  and  (not A166) );
 a48631a <=( a48630a  and  a48627a );
 a48634a <=( A203  and  A200 );
 a48637a <=( (not A235)  and  (not A234) );
 a48638a <=( a48637a  and  a48634a );
 a48639a <=( a48638a  and  a48631a );
 a48642a <=( (not A265)  and  (not A236) );
 a48645a <=( (not A268)  and  (not A266) );
 a48646a <=( a48645a  and  a48642a );
 a48649a <=( A299  and  A298 );
 a48652a <=( (not A301)  and  (not A300) );
 a48653a <=( a48652a  and  a48649a );
 a48654a <=( a48653a  and  a48646a );
 a48657a <=( (not A167)  and  (not A169) );
 a48660a <=( (not A199)  and  (not A166) );
 a48661a <=( a48660a  and  a48657a );
 a48664a <=( A203  and  A200 );
 a48667a <=( A233  and  A232 );
 a48668a <=( a48667a  and  a48664a );
 a48669a <=( a48668a  and  a48661a );
 a48672a <=( (not A235)  and  (not A234) );
 a48675a <=( (not A268)  and  (not A267) );
 a48676a <=( a48675a  and  a48672a );
 a48679a <=( (not A300)  and  (not A269) );
 a48682a <=( (not A302)  and  (not A301) );
 a48683a <=( a48682a  and  a48679a );
 a48684a <=( a48683a  and  a48676a );
 a48687a <=( (not A167)  and  (not A169) );
 a48690a <=( (not A199)  and  (not A166) );
 a48691a <=( a48690a  and  a48687a );
 a48694a <=( A203  and  A200 );
 a48697a <=( A233  and  A232 );
 a48698a <=( a48697a  and  a48694a );
 a48699a <=( a48698a  and  a48691a );
 a48702a <=( (not A235)  and  (not A234) );
 a48705a <=( (not A268)  and  (not A267) );
 a48706a <=( a48705a  and  a48702a );
 a48709a <=( (not A298)  and  (not A269) );
 a48712a <=( (not A301)  and  (not A299) );
 a48713a <=( a48712a  and  a48709a );
 a48714a <=( a48713a  and  a48706a );
 a48717a <=( (not A167)  and  (not A169) );
 a48720a <=( (not A199)  and  (not A166) );
 a48721a <=( a48720a  and  a48717a );
 a48724a <=( A203  and  A200 );
 a48727a <=( A233  and  A232 );
 a48728a <=( a48727a  and  a48724a );
 a48729a <=( a48728a  and  a48721a );
 a48732a <=( (not A235)  and  (not A234) );
 a48735a <=( (not A266)  and  (not A265) );
 a48736a <=( a48735a  and  a48732a );
 a48739a <=( (not A300)  and  (not A268) );
 a48742a <=( (not A302)  and  (not A301) );
 a48743a <=( a48742a  and  a48739a );
 a48744a <=( a48743a  and  a48736a );
 a48747a <=( (not A167)  and  (not A169) );
 a48750a <=( (not A199)  and  (not A166) );
 a48751a <=( a48750a  and  a48747a );
 a48754a <=( A203  and  A200 );
 a48757a <=( A233  and  A232 );
 a48758a <=( a48757a  and  a48754a );
 a48759a <=( a48758a  and  a48751a );
 a48762a <=( (not A235)  and  (not A234) );
 a48765a <=( (not A266)  and  (not A265) );
 a48766a <=( a48765a  and  a48762a );
 a48769a <=( (not A298)  and  (not A268) );
 a48772a <=( (not A301)  and  (not A299) );
 a48773a <=( a48772a  and  a48769a );
 a48774a <=( a48773a  and  a48766a );
 a48777a <=( (not A167)  and  (not A169) );
 a48780a <=( (not A199)  and  (not A166) );
 a48781a <=( a48780a  and  a48777a );
 a48784a <=( A203  and  A200 );
 a48787a <=( (not A233)  and  (not A232) );
 a48788a <=( a48787a  and  a48784a );
 a48789a <=( a48788a  and  a48781a );
 a48792a <=( (not A267)  and  (not A235) );
 a48795a <=( (not A269)  and  (not A268) );
 a48796a <=( a48795a  and  a48792a );
 a48799a <=( A299  and  A298 );
 a48802a <=( (not A301)  and  (not A300) );
 a48803a <=( a48802a  and  a48799a );
 a48804a <=( a48803a  and  a48796a );
 a48807a <=( (not A167)  and  (not A169) );
 a48810a <=( (not A199)  and  (not A166) );
 a48811a <=( a48810a  and  a48807a );
 a48814a <=( A203  and  A200 );
 a48817a <=( (not A233)  and  (not A232) );
 a48818a <=( a48817a  and  a48814a );
 a48819a <=( a48818a  and  a48811a );
 a48822a <=( A265  and  (not A235) );
 a48825a <=( (not A267)  and  A266 );
 a48826a <=( a48825a  and  a48822a );
 a48829a <=( (not A300)  and  (not A268) );
 a48832a <=( (not A302)  and  (not A301) );
 a48833a <=( a48832a  and  a48829a );
 a48834a <=( a48833a  and  a48826a );
 a48837a <=( (not A167)  and  (not A169) );
 a48840a <=( (not A199)  and  (not A166) );
 a48841a <=( a48840a  and  a48837a );
 a48844a <=( A203  and  A200 );
 a48847a <=( (not A233)  and  (not A232) );
 a48848a <=( a48847a  and  a48844a );
 a48849a <=( a48848a  and  a48841a );
 a48852a <=( A265  and  (not A235) );
 a48855a <=( (not A267)  and  A266 );
 a48856a <=( a48855a  and  a48852a );
 a48859a <=( (not A298)  and  (not A268) );
 a48862a <=( (not A301)  and  (not A299) );
 a48863a <=( a48862a  and  a48859a );
 a48864a <=( a48863a  and  a48856a );
 a48867a <=( (not A167)  and  (not A169) );
 a48870a <=( (not A199)  and  (not A166) );
 a48871a <=( a48870a  and  a48867a );
 a48874a <=( A203  and  A200 );
 a48877a <=( (not A233)  and  (not A232) );
 a48878a <=( a48877a  and  a48874a );
 a48879a <=( a48878a  and  a48871a );
 a48882a <=( (not A265)  and  (not A235) );
 a48885a <=( (not A268)  and  (not A266) );
 a48886a <=( a48885a  and  a48882a );
 a48889a <=( A299  and  A298 );
 a48892a <=( (not A301)  and  (not A300) );
 a48893a <=( a48892a  and  a48889a );
 a48894a <=( a48893a  and  a48886a );
 a48897a <=( (not A167)  and  (not A169) );
 a48900a <=( A199  and  (not A166) );
 a48901a <=( a48900a  and  a48897a );
 a48904a <=( A203  and  (not A200) );
 a48907a <=( (not A235)  and  (not A234) );
 a48908a <=( a48907a  and  a48904a );
 a48909a <=( a48908a  and  a48901a );
 a48912a <=( (not A267)  and  (not A236) );
 a48915a <=( (not A269)  and  (not A268) );
 a48916a <=( a48915a  and  a48912a );
 a48919a <=( A299  and  A298 );
 a48922a <=( (not A301)  and  (not A300) );
 a48923a <=( a48922a  and  a48919a );
 a48924a <=( a48923a  and  a48916a );
 a48927a <=( (not A167)  and  (not A169) );
 a48930a <=( A199  and  (not A166) );
 a48931a <=( a48930a  and  a48927a );
 a48934a <=( A203  and  (not A200) );
 a48937a <=( (not A235)  and  (not A234) );
 a48938a <=( a48937a  and  a48934a );
 a48939a <=( a48938a  and  a48931a );
 a48942a <=( A265  and  (not A236) );
 a48945a <=( (not A267)  and  A266 );
 a48946a <=( a48945a  and  a48942a );
 a48949a <=( (not A300)  and  (not A268) );
 a48952a <=( (not A302)  and  (not A301) );
 a48953a <=( a48952a  and  a48949a );
 a48954a <=( a48953a  and  a48946a );
 a48957a <=( (not A167)  and  (not A169) );
 a48960a <=( A199  and  (not A166) );
 a48961a <=( a48960a  and  a48957a );
 a48964a <=( A203  and  (not A200) );
 a48967a <=( (not A235)  and  (not A234) );
 a48968a <=( a48967a  and  a48964a );
 a48969a <=( a48968a  and  a48961a );
 a48972a <=( A265  and  (not A236) );
 a48975a <=( (not A267)  and  A266 );
 a48976a <=( a48975a  and  a48972a );
 a48979a <=( (not A298)  and  (not A268) );
 a48982a <=( (not A301)  and  (not A299) );
 a48983a <=( a48982a  and  a48979a );
 a48984a <=( a48983a  and  a48976a );
 a48987a <=( (not A167)  and  (not A169) );
 a48990a <=( A199  and  (not A166) );
 a48991a <=( a48990a  and  a48987a );
 a48994a <=( A203  and  (not A200) );
 a48997a <=( (not A235)  and  (not A234) );
 a48998a <=( a48997a  and  a48994a );
 a48999a <=( a48998a  and  a48991a );
 a49002a <=( (not A265)  and  (not A236) );
 a49005a <=( (not A268)  and  (not A266) );
 a49006a <=( a49005a  and  a49002a );
 a49009a <=( A299  and  A298 );
 a49012a <=( (not A301)  and  (not A300) );
 a49013a <=( a49012a  and  a49009a );
 a49014a <=( a49013a  and  a49006a );
 a49017a <=( (not A167)  and  (not A169) );
 a49020a <=( A199  and  (not A166) );
 a49021a <=( a49020a  and  a49017a );
 a49024a <=( A203  and  (not A200) );
 a49027a <=( A233  and  A232 );
 a49028a <=( a49027a  and  a49024a );
 a49029a <=( a49028a  and  a49021a );
 a49032a <=( (not A235)  and  (not A234) );
 a49035a <=( (not A268)  and  (not A267) );
 a49036a <=( a49035a  and  a49032a );
 a49039a <=( (not A300)  and  (not A269) );
 a49042a <=( (not A302)  and  (not A301) );
 a49043a <=( a49042a  and  a49039a );
 a49044a <=( a49043a  and  a49036a );
 a49047a <=( (not A167)  and  (not A169) );
 a49050a <=( A199  and  (not A166) );
 a49051a <=( a49050a  and  a49047a );
 a49054a <=( A203  and  (not A200) );
 a49057a <=( A233  and  A232 );
 a49058a <=( a49057a  and  a49054a );
 a49059a <=( a49058a  and  a49051a );
 a49062a <=( (not A235)  and  (not A234) );
 a49065a <=( (not A268)  and  (not A267) );
 a49066a <=( a49065a  and  a49062a );
 a49069a <=( (not A298)  and  (not A269) );
 a49072a <=( (not A301)  and  (not A299) );
 a49073a <=( a49072a  and  a49069a );
 a49074a <=( a49073a  and  a49066a );
 a49077a <=( (not A167)  and  (not A169) );
 a49080a <=( A199  and  (not A166) );
 a49081a <=( a49080a  and  a49077a );
 a49084a <=( A203  and  (not A200) );
 a49087a <=( A233  and  A232 );
 a49088a <=( a49087a  and  a49084a );
 a49089a <=( a49088a  and  a49081a );
 a49092a <=( (not A235)  and  (not A234) );
 a49095a <=( (not A266)  and  (not A265) );
 a49096a <=( a49095a  and  a49092a );
 a49099a <=( (not A300)  and  (not A268) );
 a49102a <=( (not A302)  and  (not A301) );
 a49103a <=( a49102a  and  a49099a );
 a49104a <=( a49103a  and  a49096a );
 a49107a <=( (not A167)  and  (not A169) );
 a49110a <=( A199  and  (not A166) );
 a49111a <=( a49110a  and  a49107a );
 a49114a <=( A203  and  (not A200) );
 a49117a <=( A233  and  A232 );
 a49118a <=( a49117a  and  a49114a );
 a49119a <=( a49118a  and  a49111a );
 a49122a <=( (not A235)  and  (not A234) );
 a49125a <=( (not A266)  and  (not A265) );
 a49126a <=( a49125a  and  a49122a );
 a49129a <=( (not A298)  and  (not A268) );
 a49132a <=( (not A301)  and  (not A299) );
 a49133a <=( a49132a  and  a49129a );
 a49134a <=( a49133a  and  a49126a );
 a49137a <=( (not A167)  and  (not A169) );
 a49140a <=( A199  and  (not A166) );
 a49141a <=( a49140a  and  a49137a );
 a49144a <=( A203  and  (not A200) );
 a49147a <=( (not A233)  and  (not A232) );
 a49148a <=( a49147a  and  a49144a );
 a49149a <=( a49148a  and  a49141a );
 a49152a <=( (not A267)  and  (not A235) );
 a49155a <=( (not A269)  and  (not A268) );
 a49156a <=( a49155a  and  a49152a );
 a49159a <=( A299  and  A298 );
 a49162a <=( (not A301)  and  (not A300) );
 a49163a <=( a49162a  and  a49159a );
 a49164a <=( a49163a  and  a49156a );
 a49167a <=( (not A167)  and  (not A169) );
 a49170a <=( A199  and  (not A166) );
 a49171a <=( a49170a  and  a49167a );
 a49174a <=( A203  and  (not A200) );
 a49177a <=( (not A233)  and  (not A232) );
 a49178a <=( a49177a  and  a49174a );
 a49179a <=( a49178a  and  a49171a );
 a49182a <=( A265  and  (not A235) );
 a49185a <=( (not A267)  and  A266 );
 a49186a <=( a49185a  and  a49182a );
 a49189a <=( (not A300)  and  (not A268) );
 a49192a <=( (not A302)  and  (not A301) );
 a49193a <=( a49192a  and  a49189a );
 a49194a <=( a49193a  and  a49186a );
 a49197a <=( (not A167)  and  (not A169) );
 a49200a <=( A199  and  (not A166) );
 a49201a <=( a49200a  and  a49197a );
 a49204a <=( A203  and  (not A200) );
 a49207a <=( (not A233)  and  (not A232) );
 a49208a <=( a49207a  and  a49204a );
 a49209a <=( a49208a  and  a49201a );
 a49212a <=( A265  and  (not A235) );
 a49215a <=( (not A267)  and  A266 );
 a49216a <=( a49215a  and  a49212a );
 a49219a <=( (not A298)  and  (not A268) );
 a49222a <=( (not A301)  and  (not A299) );
 a49223a <=( a49222a  and  a49219a );
 a49224a <=( a49223a  and  a49216a );
 a49227a <=( (not A167)  and  (not A169) );
 a49230a <=( A199  and  (not A166) );
 a49231a <=( a49230a  and  a49227a );
 a49234a <=( A203  and  (not A200) );
 a49237a <=( (not A233)  and  (not A232) );
 a49238a <=( a49237a  and  a49234a );
 a49239a <=( a49238a  and  a49231a );
 a49242a <=( (not A265)  and  (not A235) );
 a49245a <=( (not A268)  and  (not A266) );
 a49246a <=( a49245a  and  a49242a );
 a49249a <=( A299  and  A298 );
 a49252a <=( (not A301)  and  (not A300) );
 a49253a <=( a49252a  and  a49249a );
 a49254a <=( a49253a  and  a49246a );
 a49257a <=( (not A168)  and  (not A169) );
 a49260a <=( A166  and  A167 );
 a49261a <=( a49260a  and  a49257a );
 a49264a <=( (not A234)  and  A202 );
 a49267a <=( (not A236)  and  (not A235) );
 a49268a <=( a49267a  and  a49264a );
 a49269a <=( a49268a  and  a49261a );
 a49272a <=( A266  and  A265 );
 a49275a <=( (not A268)  and  (not A267) );
 a49276a <=( a49275a  and  a49272a );
 a49279a <=( A299  and  A298 );
 a49282a <=( (not A301)  and  (not A300) );
 a49283a <=( a49282a  and  a49279a );
 a49284a <=( a49283a  and  a49276a );
 a49287a <=( (not A168)  and  (not A169) );
 a49290a <=( A166  and  A167 );
 a49291a <=( a49290a  and  a49287a );
 a49294a <=( A232  and  A202 );
 a49297a <=( (not A234)  and  A233 );
 a49298a <=( a49297a  and  a49294a );
 a49299a <=( a49298a  and  a49291a );
 a49302a <=( (not A267)  and  (not A235) );
 a49305a <=( (not A269)  and  (not A268) );
 a49306a <=( a49305a  and  a49302a );
 a49309a <=( A299  and  A298 );
 a49312a <=( (not A301)  and  (not A300) );
 a49313a <=( a49312a  and  a49309a );
 a49314a <=( a49313a  and  a49306a );
 a49317a <=( (not A168)  and  (not A169) );
 a49320a <=( A166  and  A167 );
 a49321a <=( a49320a  and  a49317a );
 a49324a <=( A232  and  A202 );
 a49327a <=( (not A234)  and  A233 );
 a49328a <=( a49327a  and  a49324a );
 a49329a <=( a49328a  and  a49321a );
 a49332a <=( A265  and  (not A235) );
 a49335a <=( (not A267)  and  A266 );
 a49336a <=( a49335a  and  a49332a );
 a49339a <=( (not A300)  and  (not A268) );
 a49342a <=( (not A302)  and  (not A301) );
 a49343a <=( a49342a  and  a49339a );
 a49344a <=( a49343a  and  a49336a );
 a49347a <=( (not A168)  and  (not A169) );
 a49350a <=( A166  and  A167 );
 a49351a <=( a49350a  and  a49347a );
 a49354a <=( A232  and  A202 );
 a49357a <=( (not A234)  and  A233 );
 a49358a <=( a49357a  and  a49354a );
 a49359a <=( a49358a  and  a49351a );
 a49362a <=( A265  and  (not A235) );
 a49365a <=( (not A267)  and  A266 );
 a49366a <=( a49365a  and  a49362a );
 a49369a <=( (not A298)  and  (not A268) );
 a49372a <=( (not A301)  and  (not A299) );
 a49373a <=( a49372a  and  a49369a );
 a49374a <=( a49373a  and  a49366a );
 a49377a <=( (not A168)  and  (not A169) );
 a49380a <=( A166  and  A167 );
 a49381a <=( a49380a  and  a49377a );
 a49384a <=( A232  and  A202 );
 a49387a <=( (not A234)  and  A233 );
 a49388a <=( a49387a  and  a49384a );
 a49389a <=( a49388a  and  a49381a );
 a49392a <=( (not A265)  and  (not A235) );
 a49395a <=( (not A268)  and  (not A266) );
 a49396a <=( a49395a  and  a49392a );
 a49399a <=( A299  and  A298 );
 a49402a <=( (not A301)  and  (not A300) );
 a49403a <=( a49402a  and  a49399a );
 a49404a <=( a49403a  and  a49396a );
 a49407a <=( (not A168)  and  (not A169) );
 a49410a <=( A166  and  A167 );
 a49411a <=( a49410a  and  a49407a );
 a49414a <=( (not A232)  and  A202 );
 a49417a <=( (not A235)  and  (not A233) );
 a49418a <=( a49417a  and  a49414a );
 a49419a <=( a49418a  and  a49411a );
 a49422a <=( A266  and  A265 );
 a49425a <=( (not A268)  and  (not A267) );
 a49426a <=( a49425a  and  a49422a );
 a49429a <=( A299  and  A298 );
 a49432a <=( (not A301)  and  (not A300) );
 a49433a <=( a49432a  and  a49429a );
 a49434a <=( a49433a  and  a49426a );
 a49437a <=( (not A168)  and  (not A169) );
 a49440a <=( A166  and  A167 );
 a49441a <=( a49440a  and  a49437a );
 a49444a <=( A201  and  A199 );
 a49447a <=( (not A235)  and  (not A234) );
 a49448a <=( a49447a  and  a49444a );
 a49449a <=( a49448a  and  a49441a );
 a49452a <=( (not A267)  and  (not A236) );
 a49455a <=( (not A269)  and  (not A268) );
 a49456a <=( a49455a  and  a49452a );
 a49459a <=( A299  and  A298 );
 a49462a <=( (not A301)  and  (not A300) );
 a49463a <=( a49462a  and  a49459a );
 a49464a <=( a49463a  and  a49456a );
 a49467a <=( (not A168)  and  (not A169) );
 a49470a <=( A166  and  A167 );
 a49471a <=( a49470a  and  a49467a );
 a49474a <=( A201  and  A199 );
 a49477a <=( (not A235)  and  (not A234) );
 a49478a <=( a49477a  and  a49474a );
 a49479a <=( a49478a  and  a49471a );
 a49482a <=( A265  and  (not A236) );
 a49485a <=( (not A267)  and  A266 );
 a49486a <=( a49485a  and  a49482a );
 a49489a <=( (not A300)  and  (not A268) );
 a49492a <=( (not A302)  and  (not A301) );
 a49493a <=( a49492a  and  a49489a );
 a49494a <=( a49493a  and  a49486a );
 a49497a <=( (not A168)  and  (not A169) );
 a49500a <=( A166  and  A167 );
 a49501a <=( a49500a  and  a49497a );
 a49504a <=( A201  and  A199 );
 a49507a <=( (not A235)  and  (not A234) );
 a49508a <=( a49507a  and  a49504a );
 a49509a <=( a49508a  and  a49501a );
 a49512a <=( A265  and  (not A236) );
 a49515a <=( (not A267)  and  A266 );
 a49516a <=( a49515a  and  a49512a );
 a49519a <=( (not A298)  and  (not A268) );
 a49522a <=( (not A301)  and  (not A299) );
 a49523a <=( a49522a  and  a49519a );
 a49524a <=( a49523a  and  a49516a );
 a49527a <=( (not A168)  and  (not A169) );
 a49530a <=( A166  and  A167 );
 a49531a <=( a49530a  and  a49527a );
 a49534a <=( A201  and  A199 );
 a49537a <=( (not A235)  and  (not A234) );
 a49538a <=( a49537a  and  a49534a );
 a49539a <=( a49538a  and  a49531a );
 a49542a <=( (not A265)  and  (not A236) );
 a49545a <=( (not A268)  and  (not A266) );
 a49546a <=( a49545a  and  a49542a );
 a49549a <=( A299  and  A298 );
 a49552a <=( (not A301)  and  (not A300) );
 a49553a <=( a49552a  and  a49549a );
 a49554a <=( a49553a  and  a49546a );
 a49557a <=( (not A168)  and  (not A169) );
 a49560a <=( A166  and  A167 );
 a49561a <=( a49560a  and  a49557a );
 a49564a <=( A201  and  A199 );
 a49567a <=( A233  and  A232 );
 a49568a <=( a49567a  and  a49564a );
 a49569a <=( a49568a  and  a49561a );
 a49572a <=( (not A235)  and  (not A234) );
 a49575a <=( (not A268)  and  (not A267) );
 a49576a <=( a49575a  and  a49572a );
 a49579a <=( (not A300)  and  (not A269) );
 a49582a <=( (not A302)  and  (not A301) );
 a49583a <=( a49582a  and  a49579a );
 a49584a <=( a49583a  and  a49576a );
 a49587a <=( (not A168)  and  (not A169) );
 a49590a <=( A166  and  A167 );
 a49591a <=( a49590a  and  a49587a );
 a49594a <=( A201  and  A199 );
 a49597a <=( A233  and  A232 );
 a49598a <=( a49597a  and  a49594a );
 a49599a <=( a49598a  and  a49591a );
 a49602a <=( (not A235)  and  (not A234) );
 a49605a <=( (not A268)  and  (not A267) );
 a49606a <=( a49605a  and  a49602a );
 a49609a <=( (not A298)  and  (not A269) );
 a49612a <=( (not A301)  and  (not A299) );
 a49613a <=( a49612a  and  a49609a );
 a49614a <=( a49613a  and  a49606a );
 a49617a <=( (not A168)  and  (not A169) );
 a49620a <=( A166  and  A167 );
 a49621a <=( a49620a  and  a49617a );
 a49624a <=( A201  and  A199 );
 a49627a <=( A233  and  A232 );
 a49628a <=( a49627a  and  a49624a );
 a49629a <=( a49628a  and  a49621a );
 a49632a <=( (not A235)  and  (not A234) );
 a49635a <=( (not A266)  and  (not A265) );
 a49636a <=( a49635a  and  a49632a );
 a49639a <=( (not A300)  and  (not A268) );
 a49642a <=( (not A302)  and  (not A301) );
 a49643a <=( a49642a  and  a49639a );
 a49644a <=( a49643a  and  a49636a );
 a49647a <=( (not A168)  and  (not A169) );
 a49650a <=( A166  and  A167 );
 a49651a <=( a49650a  and  a49647a );
 a49654a <=( A201  and  A199 );
 a49657a <=( A233  and  A232 );
 a49658a <=( a49657a  and  a49654a );
 a49659a <=( a49658a  and  a49651a );
 a49662a <=( (not A235)  and  (not A234) );
 a49665a <=( (not A266)  and  (not A265) );
 a49666a <=( a49665a  and  a49662a );
 a49669a <=( (not A298)  and  (not A268) );
 a49672a <=( (not A301)  and  (not A299) );
 a49673a <=( a49672a  and  a49669a );
 a49674a <=( a49673a  and  a49666a );
 a49677a <=( (not A168)  and  (not A169) );
 a49680a <=( A166  and  A167 );
 a49681a <=( a49680a  and  a49677a );
 a49684a <=( A201  and  A199 );
 a49687a <=( (not A233)  and  (not A232) );
 a49688a <=( a49687a  and  a49684a );
 a49689a <=( a49688a  and  a49681a );
 a49692a <=( (not A267)  and  (not A235) );
 a49695a <=( (not A269)  and  (not A268) );
 a49696a <=( a49695a  and  a49692a );
 a49699a <=( A299  and  A298 );
 a49702a <=( (not A301)  and  (not A300) );
 a49703a <=( a49702a  and  a49699a );
 a49704a <=( a49703a  and  a49696a );
 a49707a <=( (not A168)  and  (not A169) );
 a49710a <=( A166  and  A167 );
 a49711a <=( a49710a  and  a49707a );
 a49714a <=( A201  and  A199 );
 a49717a <=( (not A233)  and  (not A232) );
 a49718a <=( a49717a  and  a49714a );
 a49719a <=( a49718a  and  a49711a );
 a49722a <=( A265  and  (not A235) );
 a49725a <=( (not A267)  and  A266 );
 a49726a <=( a49725a  and  a49722a );
 a49729a <=( (not A300)  and  (not A268) );
 a49732a <=( (not A302)  and  (not A301) );
 a49733a <=( a49732a  and  a49729a );
 a49734a <=( a49733a  and  a49726a );
 a49737a <=( (not A168)  and  (not A169) );
 a49740a <=( A166  and  A167 );
 a49741a <=( a49740a  and  a49737a );
 a49744a <=( A201  and  A199 );
 a49747a <=( (not A233)  and  (not A232) );
 a49748a <=( a49747a  and  a49744a );
 a49749a <=( a49748a  and  a49741a );
 a49752a <=( A265  and  (not A235) );
 a49755a <=( (not A267)  and  A266 );
 a49756a <=( a49755a  and  a49752a );
 a49759a <=( (not A298)  and  (not A268) );
 a49762a <=( (not A301)  and  (not A299) );
 a49763a <=( a49762a  and  a49759a );
 a49764a <=( a49763a  and  a49756a );
 a49767a <=( (not A168)  and  (not A169) );
 a49770a <=( A166  and  A167 );
 a49771a <=( a49770a  and  a49767a );
 a49774a <=( A201  and  A199 );
 a49777a <=( (not A233)  and  (not A232) );
 a49778a <=( a49777a  and  a49774a );
 a49779a <=( a49778a  and  a49771a );
 a49782a <=( (not A265)  and  (not A235) );
 a49785a <=( (not A268)  and  (not A266) );
 a49786a <=( a49785a  and  a49782a );
 a49789a <=( A299  and  A298 );
 a49792a <=( (not A301)  and  (not A300) );
 a49793a <=( a49792a  and  a49789a );
 a49794a <=( a49793a  and  a49786a );
 a49797a <=( (not A168)  and  (not A169) );
 a49800a <=( A166  and  A167 );
 a49801a <=( a49800a  and  a49797a );
 a49804a <=( A201  and  A200 );
 a49807a <=( (not A235)  and  (not A234) );
 a49808a <=( a49807a  and  a49804a );
 a49809a <=( a49808a  and  a49801a );
 a49812a <=( (not A267)  and  (not A236) );
 a49815a <=( (not A269)  and  (not A268) );
 a49816a <=( a49815a  and  a49812a );
 a49819a <=( A299  and  A298 );
 a49822a <=( (not A301)  and  (not A300) );
 a49823a <=( a49822a  and  a49819a );
 a49824a <=( a49823a  and  a49816a );
 a49827a <=( (not A168)  and  (not A169) );
 a49830a <=( A166  and  A167 );
 a49831a <=( a49830a  and  a49827a );
 a49834a <=( A201  and  A200 );
 a49837a <=( (not A235)  and  (not A234) );
 a49838a <=( a49837a  and  a49834a );
 a49839a <=( a49838a  and  a49831a );
 a49842a <=( A265  and  (not A236) );
 a49845a <=( (not A267)  and  A266 );
 a49846a <=( a49845a  and  a49842a );
 a49849a <=( (not A300)  and  (not A268) );
 a49852a <=( (not A302)  and  (not A301) );
 a49853a <=( a49852a  and  a49849a );
 a49854a <=( a49853a  and  a49846a );
 a49857a <=( (not A168)  and  (not A169) );
 a49860a <=( A166  and  A167 );
 a49861a <=( a49860a  and  a49857a );
 a49864a <=( A201  and  A200 );
 a49867a <=( (not A235)  and  (not A234) );
 a49868a <=( a49867a  and  a49864a );
 a49869a <=( a49868a  and  a49861a );
 a49872a <=( A265  and  (not A236) );
 a49875a <=( (not A267)  and  A266 );
 a49876a <=( a49875a  and  a49872a );
 a49879a <=( (not A298)  and  (not A268) );
 a49882a <=( (not A301)  and  (not A299) );
 a49883a <=( a49882a  and  a49879a );
 a49884a <=( a49883a  and  a49876a );
 a49887a <=( (not A168)  and  (not A169) );
 a49890a <=( A166  and  A167 );
 a49891a <=( a49890a  and  a49887a );
 a49894a <=( A201  and  A200 );
 a49897a <=( (not A235)  and  (not A234) );
 a49898a <=( a49897a  and  a49894a );
 a49899a <=( a49898a  and  a49891a );
 a49902a <=( (not A265)  and  (not A236) );
 a49905a <=( (not A268)  and  (not A266) );
 a49906a <=( a49905a  and  a49902a );
 a49909a <=( A299  and  A298 );
 a49912a <=( (not A301)  and  (not A300) );
 a49913a <=( a49912a  and  a49909a );
 a49914a <=( a49913a  and  a49906a );
 a49917a <=( (not A168)  and  (not A169) );
 a49920a <=( A166  and  A167 );
 a49921a <=( a49920a  and  a49917a );
 a49924a <=( A201  and  A200 );
 a49927a <=( A233  and  A232 );
 a49928a <=( a49927a  and  a49924a );
 a49929a <=( a49928a  and  a49921a );
 a49932a <=( (not A235)  and  (not A234) );
 a49935a <=( (not A268)  and  (not A267) );
 a49936a <=( a49935a  and  a49932a );
 a49939a <=( (not A300)  and  (not A269) );
 a49942a <=( (not A302)  and  (not A301) );
 a49943a <=( a49942a  and  a49939a );
 a49944a <=( a49943a  and  a49936a );
 a49947a <=( (not A168)  and  (not A169) );
 a49950a <=( A166  and  A167 );
 a49951a <=( a49950a  and  a49947a );
 a49954a <=( A201  and  A200 );
 a49957a <=( A233  and  A232 );
 a49958a <=( a49957a  and  a49954a );
 a49959a <=( a49958a  and  a49951a );
 a49962a <=( (not A235)  and  (not A234) );
 a49965a <=( (not A268)  and  (not A267) );
 a49966a <=( a49965a  and  a49962a );
 a49969a <=( (not A298)  and  (not A269) );
 a49972a <=( (not A301)  and  (not A299) );
 a49973a <=( a49972a  and  a49969a );
 a49974a <=( a49973a  and  a49966a );
 a49977a <=( (not A168)  and  (not A169) );
 a49980a <=( A166  and  A167 );
 a49981a <=( a49980a  and  a49977a );
 a49984a <=( A201  and  A200 );
 a49987a <=( A233  and  A232 );
 a49988a <=( a49987a  and  a49984a );
 a49989a <=( a49988a  and  a49981a );
 a49992a <=( (not A235)  and  (not A234) );
 a49995a <=( (not A266)  and  (not A265) );
 a49996a <=( a49995a  and  a49992a );
 a49999a <=( (not A300)  and  (not A268) );
 a50002a <=( (not A302)  and  (not A301) );
 a50003a <=( a50002a  and  a49999a );
 a50004a <=( a50003a  and  a49996a );
 a50007a <=( (not A168)  and  (not A169) );
 a50010a <=( A166  and  A167 );
 a50011a <=( a50010a  and  a50007a );
 a50014a <=( A201  and  A200 );
 a50017a <=( A233  and  A232 );
 a50018a <=( a50017a  and  a50014a );
 a50019a <=( a50018a  and  a50011a );
 a50022a <=( (not A235)  and  (not A234) );
 a50025a <=( (not A266)  and  (not A265) );
 a50026a <=( a50025a  and  a50022a );
 a50029a <=( (not A298)  and  (not A268) );
 a50032a <=( (not A301)  and  (not A299) );
 a50033a <=( a50032a  and  a50029a );
 a50034a <=( a50033a  and  a50026a );
 a50037a <=( (not A168)  and  (not A169) );
 a50040a <=( A166  and  A167 );
 a50041a <=( a50040a  and  a50037a );
 a50044a <=( A201  and  A200 );
 a50047a <=( (not A233)  and  (not A232) );
 a50048a <=( a50047a  and  a50044a );
 a50049a <=( a50048a  and  a50041a );
 a50052a <=( (not A267)  and  (not A235) );
 a50055a <=( (not A269)  and  (not A268) );
 a50056a <=( a50055a  and  a50052a );
 a50059a <=( A299  and  A298 );
 a50062a <=( (not A301)  and  (not A300) );
 a50063a <=( a50062a  and  a50059a );
 a50064a <=( a50063a  and  a50056a );
 a50067a <=( (not A168)  and  (not A169) );
 a50070a <=( A166  and  A167 );
 a50071a <=( a50070a  and  a50067a );
 a50074a <=( A201  and  A200 );
 a50077a <=( (not A233)  and  (not A232) );
 a50078a <=( a50077a  and  a50074a );
 a50079a <=( a50078a  and  a50071a );
 a50082a <=( A265  and  (not A235) );
 a50085a <=( (not A267)  and  A266 );
 a50086a <=( a50085a  and  a50082a );
 a50089a <=( (not A300)  and  (not A268) );
 a50092a <=( (not A302)  and  (not A301) );
 a50093a <=( a50092a  and  a50089a );
 a50094a <=( a50093a  and  a50086a );
 a50097a <=( (not A168)  and  (not A169) );
 a50100a <=( A166  and  A167 );
 a50101a <=( a50100a  and  a50097a );
 a50104a <=( A201  and  A200 );
 a50107a <=( (not A233)  and  (not A232) );
 a50108a <=( a50107a  and  a50104a );
 a50109a <=( a50108a  and  a50101a );
 a50112a <=( A265  and  (not A235) );
 a50115a <=( (not A267)  and  A266 );
 a50116a <=( a50115a  and  a50112a );
 a50119a <=( (not A298)  and  (not A268) );
 a50122a <=( (not A301)  and  (not A299) );
 a50123a <=( a50122a  and  a50119a );
 a50124a <=( a50123a  and  a50116a );
 a50127a <=( (not A168)  and  (not A169) );
 a50130a <=( A166  and  A167 );
 a50131a <=( a50130a  and  a50127a );
 a50134a <=( A201  and  A200 );
 a50137a <=( (not A233)  and  (not A232) );
 a50138a <=( a50137a  and  a50134a );
 a50139a <=( a50138a  and  a50131a );
 a50142a <=( (not A265)  and  (not A235) );
 a50145a <=( (not A268)  and  (not A266) );
 a50146a <=( a50145a  and  a50142a );
 a50149a <=( A299  and  A298 );
 a50152a <=( (not A301)  and  (not A300) );
 a50153a <=( a50152a  and  a50149a );
 a50154a <=( a50153a  and  a50146a );
 a50157a <=( (not A168)  and  (not A169) );
 a50160a <=( A166  and  A167 );
 a50161a <=( a50160a  and  a50157a );
 a50164a <=( A200  and  (not A199) );
 a50167a <=( (not A234)  and  A203 );
 a50168a <=( a50167a  and  a50164a );
 a50169a <=( a50168a  and  a50161a );
 a50172a <=( (not A236)  and  (not A235) );
 a50175a <=( (not A268)  and  (not A267) );
 a50176a <=( a50175a  and  a50172a );
 a50179a <=( (not A300)  and  (not A269) );
 a50182a <=( (not A302)  and  (not A301) );
 a50183a <=( a50182a  and  a50179a );
 a50184a <=( a50183a  and  a50176a );
 a50187a <=( (not A168)  and  (not A169) );
 a50190a <=( A166  and  A167 );
 a50191a <=( a50190a  and  a50187a );
 a50194a <=( A200  and  (not A199) );
 a50197a <=( (not A234)  and  A203 );
 a50198a <=( a50197a  and  a50194a );
 a50199a <=( a50198a  and  a50191a );
 a50202a <=( (not A236)  and  (not A235) );
 a50205a <=( (not A268)  and  (not A267) );
 a50206a <=( a50205a  and  a50202a );
 a50209a <=( (not A298)  and  (not A269) );
 a50212a <=( (not A301)  and  (not A299) );
 a50213a <=( a50212a  and  a50209a );
 a50214a <=( a50213a  and  a50206a );
 a50217a <=( (not A168)  and  (not A169) );
 a50220a <=( A166  and  A167 );
 a50221a <=( a50220a  and  a50217a );
 a50224a <=( A200  and  (not A199) );
 a50227a <=( (not A234)  and  A203 );
 a50228a <=( a50227a  and  a50224a );
 a50229a <=( a50228a  and  a50221a );
 a50232a <=( (not A236)  and  (not A235) );
 a50235a <=( (not A266)  and  (not A265) );
 a50236a <=( a50235a  and  a50232a );
 a50239a <=( (not A300)  and  (not A268) );
 a50242a <=( (not A302)  and  (not A301) );
 a50243a <=( a50242a  and  a50239a );
 a50244a <=( a50243a  and  a50236a );
 a50247a <=( (not A168)  and  (not A169) );
 a50250a <=( A166  and  A167 );
 a50251a <=( a50250a  and  a50247a );
 a50254a <=( A200  and  (not A199) );
 a50257a <=( (not A234)  and  A203 );
 a50258a <=( a50257a  and  a50254a );
 a50259a <=( a50258a  and  a50251a );
 a50262a <=( (not A236)  and  (not A235) );
 a50265a <=( (not A266)  and  (not A265) );
 a50266a <=( a50265a  and  a50262a );
 a50269a <=( (not A298)  and  (not A268) );
 a50272a <=( (not A301)  and  (not A299) );
 a50273a <=( a50272a  and  a50269a );
 a50274a <=( a50273a  and  a50266a );
 a50277a <=( (not A168)  and  (not A169) );
 a50280a <=( A166  and  A167 );
 a50281a <=( a50280a  and  a50277a );
 a50284a <=( A200  and  (not A199) );
 a50287a <=( (not A232)  and  A203 );
 a50288a <=( a50287a  and  a50284a );
 a50289a <=( a50288a  and  a50281a );
 a50292a <=( (not A235)  and  (not A233) );
 a50295a <=( (not A268)  and  (not A267) );
 a50296a <=( a50295a  and  a50292a );
 a50299a <=( (not A300)  and  (not A269) );
 a50302a <=( (not A302)  and  (not A301) );
 a50303a <=( a50302a  and  a50299a );
 a50304a <=( a50303a  and  a50296a );
 a50307a <=( (not A168)  and  (not A169) );
 a50310a <=( A166  and  A167 );
 a50311a <=( a50310a  and  a50307a );
 a50314a <=( A200  and  (not A199) );
 a50317a <=( (not A232)  and  A203 );
 a50318a <=( a50317a  and  a50314a );
 a50319a <=( a50318a  and  a50311a );
 a50322a <=( (not A235)  and  (not A233) );
 a50325a <=( (not A268)  and  (not A267) );
 a50326a <=( a50325a  and  a50322a );
 a50329a <=( (not A298)  and  (not A269) );
 a50332a <=( (not A301)  and  (not A299) );
 a50333a <=( a50332a  and  a50329a );
 a50334a <=( a50333a  and  a50326a );
 a50337a <=( (not A168)  and  (not A169) );
 a50340a <=( A166  and  A167 );
 a50341a <=( a50340a  and  a50337a );
 a50344a <=( A200  and  (not A199) );
 a50347a <=( (not A232)  and  A203 );
 a50348a <=( a50347a  and  a50344a );
 a50349a <=( a50348a  and  a50341a );
 a50352a <=( (not A235)  and  (not A233) );
 a50355a <=( (not A266)  and  (not A265) );
 a50356a <=( a50355a  and  a50352a );
 a50359a <=( (not A300)  and  (not A268) );
 a50362a <=( (not A302)  and  (not A301) );
 a50363a <=( a50362a  and  a50359a );
 a50364a <=( a50363a  and  a50356a );
 a50367a <=( (not A168)  and  (not A169) );
 a50370a <=( A166  and  A167 );
 a50371a <=( a50370a  and  a50367a );
 a50374a <=( A200  and  (not A199) );
 a50377a <=( (not A232)  and  A203 );
 a50378a <=( a50377a  and  a50374a );
 a50379a <=( a50378a  and  a50371a );
 a50382a <=( (not A235)  and  (not A233) );
 a50385a <=( (not A266)  and  (not A265) );
 a50386a <=( a50385a  and  a50382a );
 a50389a <=( (not A298)  and  (not A268) );
 a50392a <=( (not A301)  and  (not A299) );
 a50393a <=( a50392a  and  a50389a );
 a50394a <=( a50393a  and  a50386a );
 a50397a <=( (not A168)  and  (not A169) );
 a50400a <=( A166  and  A167 );
 a50401a <=( a50400a  and  a50397a );
 a50404a <=( (not A200)  and  A199 );
 a50407a <=( (not A234)  and  A203 );
 a50408a <=( a50407a  and  a50404a );
 a50409a <=( a50408a  and  a50401a );
 a50412a <=( (not A236)  and  (not A235) );
 a50415a <=( (not A268)  and  (not A267) );
 a50416a <=( a50415a  and  a50412a );
 a50419a <=( (not A300)  and  (not A269) );
 a50422a <=( (not A302)  and  (not A301) );
 a50423a <=( a50422a  and  a50419a );
 a50424a <=( a50423a  and  a50416a );
 a50427a <=( (not A168)  and  (not A169) );
 a50430a <=( A166  and  A167 );
 a50431a <=( a50430a  and  a50427a );
 a50434a <=( (not A200)  and  A199 );
 a50437a <=( (not A234)  and  A203 );
 a50438a <=( a50437a  and  a50434a );
 a50439a <=( a50438a  and  a50431a );
 a50442a <=( (not A236)  and  (not A235) );
 a50445a <=( (not A268)  and  (not A267) );
 a50446a <=( a50445a  and  a50442a );
 a50449a <=( (not A298)  and  (not A269) );
 a50452a <=( (not A301)  and  (not A299) );
 a50453a <=( a50452a  and  a50449a );
 a50454a <=( a50453a  and  a50446a );
 a50457a <=( (not A168)  and  (not A169) );
 a50460a <=( A166  and  A167 );
 a50461a <=( a50460a  and  a50457a );
 a50464a <=( (not A200)  and  A199 );
 a50467a <=( (not A234)  and  A203 );
 a50468a <=( a50467a  and  a50464a );
 a50469a <=( a50468a  and  a50461a );
 a50472a <=( (not A236)  and  (not A235) );
 a50475a <=( (not A266)  and  (not A265) );
 a50476a <=( a50475a  and  a50472a );
 a50479a <=( (not A300)  and  (not A268) );
 a50482a <=( (not A302)  and  (not A301) );
 a50483a <=( a50482a  and  a50479a );
 a50484a <=( a50483a  and  a50476a );
 a50487a <=( (not A168)  and  (not A169) );
 a50490a <=( A166  and  A167 );
 a50491a <=( a50490a  and  a50487a );
 a50494a <=( (not A200)  and  A199 );
 a50497a <=( (not A234)  and  A203 );
 a50498a <=( a50497a  and  a50494a );
 a50499a <=( a50498a  and  a50491a );
 a50502a <=( (not A236)  and  (not A235) );
 a50505a <=( (not A266)  and  (not A265) );
 a50506a <=( a50505a  and  a50502a );
 a50509a <=( (not A298)  and  (not A268) );
 a50512a <=( (not A301)  and  (not A299) );
 a50513a <=( a50512a  and  a50509a );
 a50514a <=( a50513a  and  a50506a );
 a50517a <=( (not A168)  and  (not A169) );
 a50520a <=( A166  and  A167 );
 a50521a <=( a50520a  and  a50517a );
 a50524a <=( (not A200)  and  A199 );
 a50527a <=( (not A232)  and  A203 );
 a50528a <=( a50527a  and  a50524a );
 a50529a <=( a50528a  and  a50521a );
 a50532a <=( (not A235)  and  (not A233) );
 a50535a <=( (not A268)  and  (not A267) );
 a50536a <=( a50535a  and  a50532a );
 a50539a <=( (not A300)  and  (not A269) );
 a50542a <=( (not A302)  and  (not A301) );
 a50543a <=( a50542a  and  a50539a );
 a50544a <=( a50543a  and  a50536a );
 a50547a <=( (not A168)  and  (not A169) );
 a50550a <=( A166  and  A167 );
 a50551a <=( a50550a  and  a50547a );
 a50554a <=( (not A200)  and  A199 );
 a50557a <=( (not A232)  and  A203 );
 a50558a <=( a50557a  and  a50554a );
 a50559a <=( a50558a  and  a50551a );
 a50562a <=( (not A235)  and  (not A233) );
 a50565a <=( (not A268)  and  (not A267) );
 a50566a <=( a50565a  and  a50562a );
 a50569a <=( (not A298)  and  (not A269) );
 a50572a <=( (not A301)  and  (not A299) );
 a50573a <=( a50572a  and  a50569a );
 a50574a <=( a50573a  and  a50566a );
 a50577a <=( (not A168)  and  (not A169) );
 a50580a <=( A166  and  A167 );
 a50581a <=( a50580a  and  a50577a );
 a50584a <=( (not A200)  and  A199 );
 a50587a <=( (not A232)  and  A203 );
 a50588a <=( a50587a  and  a50584a );
 a50589a <=( a50588a  and  a50581a );
 a50592a <=( (not A235)  and  (not A233) );
 a50595a <=( (not A266)  and  (not A265) );
 a50596a <=( a50595a  and  a50592a );
 a50599a <=( (not A300)  and  (not A268) );
 a50602a <=( (not A302)  and  (not A301) );
 a50603a <=( a50602a  and  a50599a );
 a50604a <=( a50603a  and  a50596a );
 a50607a <=( (not A168)  and  (not A169) );
 a50610a <=( A166  and  A167 );
 a50611a <=( a50610a  and  a50607a );
 a50614a <=( (not A200)  and  A199 );
 a50617a <=( (not A232)  and  A203 );
 a50618a <=( a50617a  and  a50614a );
 a50619a <=( a50618a  and  a50611a );
 a50622a <=( (not A235)  and  (not A233) );
 a50625a <=( (not A266)  and  (not A265) );
 a50626a <=( a50625a  and  a50622a );
 a50629a <=( (not A298)  and  (not A268) );
 a50632a <=( (not A301)  and  (not A299) );
 a50633a <=( a50632a  and  a50629a );
 a50634a <=( a50633a  and  a50626a );
 a50637a <=( (not A169)  and  (not A170) );
 a50640a <=( A202  and  (not A168) );
 a50641a <=( a50640a  and  a50637a );
 a50644a <=( A233  and  A232 );
 a50647a <=( (not A235)  and  (not A234) );
 a50648a <=( a50647a  and  a50644a );
 a50649a <=( a50648a  and  a50641a );
 a50652a <=( A266  and  A265 );
 a50655a <=( (not A268)  and  (not A267) );
 a50656a <=( a50655a  and  a50652a );
 a50659a <=( A299  and  A298 );
 a50662a <=( (not A301)  and  (not A300) );
 a50663a <=( a50662a  and  a50659a );
 a50664a <=( a50663a  and  a50656a );
 a50667a <=( (not A169)  and  (not A170) );
 a50670a <=( A199  and  (not A168) );
 a50671a <=( a50670a  and  a50667a );
 a50674a <=( (not A234)  and  A201 );
 a50677a <=( (not A236)  and  (not A235) );
 a50678a <=( a50677a  and  a50674a );
 a50679a <=( a50678a  and  a50671a );
 a50682a <=( A266  and  A265 );
 a50685a <=( (not A268)  and  (not A267) );
 a50686a <=( a50685a  and  a50682a );
 a50689a <=( A299  and  A298 );
 a50692a <=( (not A301)  and  (not A300) );
 a50693a <=( a50692a  and  a50689a );
 a50694a <=( a50693a  and  a50686a );
 a50697a <=( (not A169)  and  (not A170) );
 a50700a <=( A199  and  (not A168) );
 a50701a <=( a50700a  and  a50697a );
 a50704a <=( A232  and  A201 );
 a50707a <=( (not A234)  and  A233 );
 a50708a <=( a50707a  and  a50704a );
 a50709a <=( a50708a  and  a50701a );
 a50712a <=( (not A267)  and  (not A235) );
 a50715a <=( (not A269)  and  (not A268) );
 a50716a <=( a50715a  and  a50712a );
 a50719a <=( A299  and  A298 );
 a50722a <=( (not A301)  and  (not A300) );
 a50723a <=( a50722a  and  a50719a );
 a50724a <=( a50723a  and  a50716a );
 a50727a <=( (not A169)  and  (not A170) );
 a50730a <=( A199  and  (not A168) );
 a50731a <=( a50730a  and  a50727a );
 a50734a <=( A232  and  A201 );
 a50737a <=( (not A234)  and  A233 );
 a50738a <=( a50737a  and  a50734a );
 a50739a <=( a50738a  and  a50731a );
 a50742a <=( A265  and  (not A235) );
 a50745a <=( (not A267)  and  A266 );
 a50746a <=( a50745a  and  a50742a );
 a50749a <=( (not A300)  and  (not A268) );
 a50752a <=( (not A302)  and  (not A301) );
 a50753a <=( a50752a  and  a50749a );
 a50754a <=( a50753a  and  a50746a );
 a50757a <=( (not A169)  and  (not A170) );
 a50760a <=( A199  and  (not A168) );
 a50761a <=( a50760a  and  a50757a );
 a50764a <=( A232  and  A201 );
 a50767a <=( (not A234)  and  A233 );
 a50768a <=( a50767a  and  a50764a );
 a50769a <=( a50768a  and  a50761a );
 a50772a <=( A265  and  (not A235) );
 a50775a <=( (not A267)  and  A266 );
 a50776a <=( a50775a  and  a50772a );
 a50779a <=( (not A298)  and  (not A268) );
 a50782a <=( (not A301)  and  (not A299) );
 a50783a <=( a50782a  and  a50779a );
 a50784a <=( a50783a  and  a50776a );
 a50787a <=( (not A169)  and  (not A170) );
 a50790a <=( A199  and  (not A168) );
 a50791a <=( a50790a  and  a50787a );
 a50794a <=( A232  and  A201 );
 a50797a <=( (not A234)  and  A233 );
 a50798a <=( a50797a  and  a50794a );
 a50799a <=( a50798a  and  a50791a );
 a50802a <=( (not A265)  and  (not A235) );
 a50805a <=( (not A268)  and  (not A266) );
 a50806a <=( a50805a  and  a50802a );
 a50809a <=( A299  and  A298 );
 a50812a <=( (not A301)  and  (not A300) );
 a50813a <=( a50812a  and  a50809a );
 a50814a <=( a50813a  and  a50806a );
 a50817a <=( (not A169)  and  (not A170) );
 a50820a <=( A199  and  (not A168) );
 a50821a <=( a50820a  and  a50817a );
 a50824a <=( (not A232)  and  A201 );
 a50827a <=( (not A235)  and  (not A233) );
 a50828a <=( a50827a  and  a50824a );
 a50829a <=( a50828a  and  a50821a );
 a50832a <=( A266  and  A265 );
 a50835a <=( (not A268)  and  (not A267) );
 a50836a <=( a50835a  and  a50832a );
 a50839a <=( A299  and  A298 );
 a50842a <=( (not A301)  and  (not A300) );
 a50843a <=( a50842a  and  a50839a );
 a50844a <=( a50843a  and  a50836a );
 a50847a <=( (not A169)  and  (not A170) );
 a50850a <=( A200  and  (not A168) );
 a50851a <=( a50850a  and  a50847a );
 a50854a <=( (not A234)  and  A201 );
 a50857a <=( (not A236)  and  (not A235) );
 a50858a <=( a50857a  and  a50854a );
 a50859a <=( a50858a  and  a50851a );
 a50862a <=( A266  and  A265 );
 a50865a <=( (not A268)  and  (not A267) );
 a50866a <=( a50865a  and  a50862a );
 a50869a <=( A299  and  A298 );
 a50872a <=( (not A301)  and  (not A300) );
 a50873a <=( a50872a  and  a50869a );
 a50874a <=( a50873a  and  a50866a );
 a50877a <=( (not A169)  and  (not A170) );
 a50880a <=( A200  and  (not A168) );
 a50881a <=( a50880a  and  a50877a );
 a50884a <=( A232  and  A201 );
 a50887a <=( (not A234)  and  A233 );
 a50888a <=( a50887a  and  a50884a );
 a50889a <=( a50888a  and  a50881a );
 a50892a <=( (not A267)  and  (not A235) );
 a50895a <=( (not A269)  and  (not A268) );
 a50896a <=( a50895a  and  a50892a );
 a50899a <=( A299  and  A298 );
 a50902a <=( (not A301)  and  (not A300) );
 a50903a <=( a50902a  and  a50899a );
 a50904a <=( a50903a  and  a50896a );
 a50907a <=( (not A169)  and  (not A170) );
 a50910a <=( A200  and  (not A168) );
 a50911a <=( a50910a  and  a50907a );
 a50914a <=( A232  and  A201 );
 a50917a <=( (not A234)  and  A233 );
 a50918a <=( a50917a  and  a50914a );
 a50919a <=( a50918a  and  a50911a );
 a50922a <=( A265  and  (not A235) );
 a50925a <=( (not A267)  and  A266 );
 a50926a <=( a50925a  and  a50922a );
 a50929a <=( (not A300)  and  (not A268) );
 a50932a <=( (not A302)  and  (not A301) );
 a50933a <=( a50932a  and  a50929a );
 a50934a <=( a50933a  and  a50926a );
 a50937a <=( (not A169)  and  (not A170) );
 a50940a <=( A200  and  (not A168) );
 a50941a <=( a50940a  and  a50937a );
 a50944a <=( A232  and  A201 );
 a50947a <=( (not A234)  and  A233 );
 a50948a <=( a50947a  and  a50944a );
 a50949a <=( a50948a  and  a50941a );
 a50952a <=( A265  and  (not A235) );
 a50955a <=( (not A267)  and  A266 );
 a50956a <=( a50955a  and  a50952a );
 a50959a <=( (not A298)  and  (not A268) );
 a50962a <=( (not A301)  and  (not A299) );
 a50963a <=( a50962a  and  a50959a );
 a50964a <=( a50963a  and  a50956a );
 a50967a <=( (not A169)  and  (not A170) );
 a50970a <=( A200  and  (not A168) );
 a50971a <=( a50970a  and  a50967a );
 a50974a <=( A232  and  A201 );
 a50977a <=( (not A234)  and  A233 );
 a50978a <=( a50977a  and  a50974a );
 a50979a <=( a50978a  and  a50971a );
 a50982a <=( (not A265)  and  (not A235) );
 a50985a <=( (not A268)  and  (not A266) );
 a50986a <=( a50985a  and  a50982a );
 a50989a <=( A299  and  A298 );
 a50992a <=( (not A301)  and  (not A300) );
 a50993a <=( a50992a  and  a50989a );
 a50994a <=( a50993a  and  a50986a );
 a50997a <=( (not A169)  and  (not A170) );
 a51000a <=( A200  and  (not A168) );
 a51001a <=( a51000a  and  a50997a );
 a51004a <=( (not A232)  and  A201 );
 a51007a <=( (not A235)  and  (not A233) );
 a51008a <=( a51007a  and  a51004a );
 a51009a <=( a51008a  and  a51001a );
 a51012a <=( A266  and  A265 );
 a51015a <=( (not A268)  and  (not A267) );
 a51016a <=( a51015a  and  a51012a );
 a51019a <=( A299  and  A298 );
 a51022a <=( (not A301)  and  (not A300) );
 a51023a <=( a51022a  and  a51019a );
 a51024a <=( a51023a  and  a51016a );
 a51027a <=( (not A169)  and  (not A170) );
 a51030a <=( (not A199)  and  (not A168) );
 a51031a <=( a51030a  and  a51027a );
 a51034a <=( A203  and  A200 );
 a51037a <=( (not A235)  and  (not A234) );
 a51038a <=( a51037a  and  a51034a );
 a51039a <=( a51038a  and  a51031a );
 a51042a <=( (not A267)  and  (not A236) );
 a51045a <=( (not A269)  and  (not A268) );
 a51046a <=( a51045a  and  a51042a );
 a51049a <=( A299  and  A298 );
 a51052a <=( (not A301)  and  (not A300) );
 a51053a <=( a51052a  and  a51049a );
 a51054a <=( a51053a  and  a51046a );
 a51057a <=( (not A169)  and  (not A170) );
 a51060a <=( (not A199)  and  (not A168) );
 a51061a <=( a51060a  and  a51057a );
 a51064a <=( A203  and  A200 );
 a51067a <=( (not A235)  and  (not A234) );
 a51068a <=( a51067a  and  a51064a );
 a51069a <=( a51068a  and  a51061a );
 a51072a <=( A265  and  (not A236) );
 a51075a <=( (not A267)  and  A266 );
 a51076a <=( a51075a  and  a51072a );
 a51079a <=( (not A300)  and  (not A268) );
 a51082a <=( (not A302)  and  (not A301) );
 a51083a <=( a51082a  and  a51079a );
 a51084a <=( a51083a  and  a51076a );
 a51087a <=( (not A169)  and  (not A170) );
 a51090a <=( (not A199)  and  (not A168) );
 a51091a <=( a51090a  and  a51087a );
 a51094a <=( A203  and  A200 );
 a51097a <=( (not A235)  and  (not A234) );
 a51098a <=( a51097a  and  a51094a );
 a51099a <=( a51098a  and  a51091a );
 a51102a <=( A265  and  (not A236) );
 a51105a <=( (not A267)  and  A266 );
 a51106a <=( a51105a  and  a51102a );
 a51109a <=( (not A298)  and  (not A268) );
 a51112a <=( (not A301)  and  (not A299) );
 a51113a <=( a51112a  and  a51109a );
 a51114a <=( a51113a  and  a51106a );
 a51117a <=( (not A169)  and  (not A170) );
 a51120a <=( (not A199)  and  (not A168) );
 a51121a <=( a51120a  and  a51117a );
 a51124a <=( A203  and  A200 );
 a51127a <=( (not A235)  and  (not A234) );
 a51128a <=( a51127a  and  a51124a );
 a51129a <=( a51128a  and  a51121a );
 a51132a <=( (not A265)  and  (not A236) );
 a51135a <=( (not A268)  and  (not A266) );
 a51136a <=( a51135a  and  a51132a );
 a51139a <=( A299  and  A298 );
 a51142a <=( (not A301)  and  (not A300) );
 a51143a <=( a51142a  and  a51139a );
 a51144a <=( a51143a  and  a51136a );
 a51147a <=( (not A169)  and  (not A170) );
 a51150a <=( (not A199)  and  (not A168) );
 a51151a <=( a51150a  and  a51147a );
 a51154a <=( A203  and  A200 );
 a51157a <=( A233  and  A232 );
 a51158a <=( a51157a  and  a51154a );
 a51159a <=( a51158a  and  a51151a );
 a51162a <=( (not A235)  and  (not A234) );
 a51165a <=( (not A268)  and  (not A267) );
 a51166a <=( a51165a  and  a51162a );
 a51169a <=( (not A300)  and  (not A269) );
 a51172a <=( (not A302)  and  (not A301) );
 a51173a <=( a51172a  and  a51169a );
 a51174a <=( a51173a  and  a51166a );
 a51177a <=( (not A169)  and  (not A170) );
 a51180a <=( (not A199)  and  (not A168) );
 a51181a <=( a51180a  and  a51177a );
 a51184a <=( A203  and  A200 );
 a51187a <=( A233  and  A232 );
 a51188a <=( a51187a  and  a51184a );
 a51189a <=( a51188a  and  a51181a );
 a51192a <=( (not A235)  and  (not A234) );
 a51195a <=( (not A268)  and  (not A267) );
 a51196a <=( a51195a  and  a51192a );
 a51199a <=( (not A298)  and  (not A269) );
 a51202a <=( (not A301)  and  (not A299) );
 a51203a <=( a51202a  and  a51199a );
 a51204a <=( a51203a  and  a51196a );
 a51207a <=( (not A169)  and  (not A170) );
 a51210a <=( (not A199)  and  (not A168) );
 a51211a <=( a51210a  and  a51207a );
 a51214a <=( A203  and  A200 );
 a51217a <=( A233  and  A232 );
 a51218a <=( a51217a  and  a51214a );
 a51219a <=( a51218a  and  a51211a );
 a51222a <=( (not A235)  and  (not A234) );
 a51225a <=( (not A266)  and  (not A265) );
 a51226a <=( a51225a  and  a51222a );
 a51229a <=( (not A300)  and  (not A268) );
 a51232a <=( (not A302)  and  (not A301) );
 a51233a <=( a51232a  and  a51229a );
 a51234a <=( a51233a  and  a51226a );
 a51237a <=( (not A169)  and  (not A170) );
 a51240a <=( (not A199)  and  (not A168) );
 a51241a <=( a51240a  and  a51237a );
 a51244a <=( A203  and  A200 );
 a51247a <=( A233  and  A232 );
 a51248a <=( a51247a  and  a51244a );
 a51249a <=( a51248a  and  a51241a );
 a51252a <=( (not A235)  and  (not A234) );
 a51255a <=( (not A266)  and  (not A265) );
 a51256a <=( a51255a  and  a51252a );
 a51259a <=( (not A298)  and  (not A268) );
 a51262a <=( (not A301)  and  (not A299) );
 a51263a <=( a51262a  and  a51259a );
 a51264a <=( a51263a  and  a51256a );
 a51267a <=( (not A169)  and  (not A170) );
 a51270a <=( (not A199)  and  (not A168) );
 a51271a <=( a51270a  and  a51267a );
 a51274a <=( A203  and  A200 );
 a51277a <=( (not A233)  and  (not A232) );
 a51278a <=( a51277a  and  a51274a );
 a51279a <=( a51278a  and  a51271a );
 a51282a <=( (not A267)  and  (not A235) );
 a51285a <=( (not A269)  and  (not A268) );
 a51286a <=( a51285a  and  a51282a );
 a51289a <=( A299  and  A298 );
 a51292a <=( (not A301)  and  (not A300) );
 a51293a <=( a51292a  and  a51289a );
 a51294a <=( a51293a  and  a51286a );
 a51297a <=( (not A169)  and  (not A170) );
 a51300a <=( (not A199)  and  (not A168) );
 a51301a <=( a51300a  and  a51297a );
 a51304a <=( A203  and  A200 );
 a51307a <=( (not A233)  and  (not A232) );
 a51308a <=( a51307a  and  a51304a );
 a51309a <=( a51308a  and  a51301a );
 a51312a <=( A265  and  (not A235) );
 a51315a <=( (not A267)  and  A266 );
 a51316a <=( a51315a  and  a51312a );
 a51319a <=( (not A300)  and  (not A268) );
 a51322a <=( (not A302)  and  (not A301) );
 a51323a <=( a51322a  and  a51319a );
 a51324a <=( a51323a  and  a51316a );
 a51327a <=( (not A169)  and  (not A170) );
 a51330a <=( (not A199)  and  (not A168) );
 a51331a <=( a51330a  and  a51327a );
 a51334a <=( A203  and  A200 );
 a51337a <=( (not A233)  and  (not A232) );
 a51338a <=( a51337a  and  a51334a );
 a51339a <=( a51338a  and  a51331a );
 a51342a <=( A265  and  (not A235) );
 a51345a <=( (not A267)  and  A266 );
 a51346a <=( a51345a  and  a51342a );
 a51349a <=( (not A298)  and  (not A268) );
 a51352a <=( (not A301)  and  (not A299) );
 a51353a <=( a51352a  and  a51349a );
 a51354a <=( a51353a  and  a51346a );
 a51357a <=( (not A169)  and  (not A170) );
 a51360a <=( (not A199)  and  (not A168) );
 a51361a <=( a51360a  and  a51357a );
 a51364a <=( A203  and  A200 );
 a51367a <=( (not A233)  and  (not A232) );
 a51368a <=( a51367a  and  a51364a );
 a51369a <=( a51368a  and  a51361a );
 a51372a <=( (not A265)  and  (not A235) );
 a51375a <=( (not A268)  and  (not A266) );
 a51376a <=( a51375a  and  a51372a );
 a51379a <=( A299  and  A298 );
 a51382a <=( (not A301)  and  (not A300) );
 a51383a <=( a51382a  and  a51379a );
 a51384a <=( a51383a  and  a51376a );
 a51387a <=( (not A169)  and  (not A170) );
 a51390a <=( A199  and  (not A168) );
 a51391a <=( a51390a  and  a51387a );
 a51394a <=( A203  and  (not A200) );
 a51397a <=( (not A235)  and  (not A234) );
 a51398a <=( a51397a  and  a51394a );
 a51399a <=( a51398a  and  a51391a );
 a51402a <=( (not A267)  and  (not A236) );
 a51405a <=( (not A269)  and  (not A268) );
 a51406a <=( a51405a  and  a51402a );
 a51409a <=( A299  and  A298 );
 a51412a <=( (not A301)  and  (not A300) );
 a51413a <=( a51412a  and  a51409a );
 a51414a <=( a51413a  and  a51406a );
 a51417a <=( (not A169)  and  (not A170) );
 a51420a <=( A199  and  (not A168) );
 a51421a <=( a51420a  and  a51417a );
 a51424a <=( A203  and  (not A200) );
 a51427a <=( (not A235)  and  (not A234) );
 a51428a <=( a51427a  and  a51424a );
 a51429a <=( a51428a  and  a51421a );
 a51432a <=( A265  and  (not A236) );
 a51435a <=( (not A267)  and  A266 );
 a51436a <=( a51435a  and  a51432a );
 a51439a <=( (not A300)  and  (not A268) );
 a51442a <=( (not A302)  and  (not A301) );
 a51443a <=( a51442a  and  a51439a );
 a51444a <=( a51443a  and  a51436a );
 a51447a <=( (not A169)  and  (not A170) );
 a51450a <=( A199  and  (not A168) );
 a51451a <=( a51450a  and  a51447a );
 a51454a <=( A203  and  (not A200) );
 a51457a <=( (not A235)  and  (not A234) );
 a51458a <=( a51457a  and  a51454a );
 a51459a <=( a51458a  and  a51451a );
 a51462a <=( A265  and  (not A236) );
 a51465a <=( (not A267)  and  A266 );
 a51466a <=( a51465a  and  a51462a );
 a51469a <=( (not A298)  and  (not A268) );
 a51472a <=( (not A301)  and  (not A299) );
 a51473a <=( a51472a  and  a51469a );
 a51474a <=( a51473a  and  a51466a );
 a51477a <=( (not A169)  and  (not A170) );
 a51480a <=( A199  and  (not A168) );
 a51481a <=( a51480a  and  a51477a );
 a51484a <=( A203  and  (not A200) );
 a51487a <=( (not A235)  and  (not A234) );
 a51488a <=( a51487a  and  a51484a );
 a51489a <=( a51488a  and  a51481a );
 a51492a <=( (not A265)  and  (not A236) );
 a51495a <=( (not A268)  and  (not A266) );
 a51496a <=( a51495a  and  a51492a );
 a51499a <=( A299  and  A298 );
 a51502a <=( (not A301)  and  (not A300) );
 a51503a <=( a51502a  and  a51499a );
 a51504a <=( a51503a  and  a51496a );
 a51507a <=( (not A169)  and  (not A170) );
 a51510a <=( A199  and  (not A168) );
 a51511a <=( a51510a  and  a51507a );
 a51514a <=( A203  and  (not A200) );
 a51517a <=( A233  and  A232 );
 a51518a <=( a51517a  and  a51514a );
 a51519a <=( a51518a  and  a51511a );
 a51522a <=( (not A235)  and  (not A234) );
 a51525a <=( (not A268)  and  (not A267) );
 a51526a <=( a51525a  and  a51522a );
 a51529a <=( (not A300)  and  (not A269) );
 a51532a <=( (not A302)  and  (not A301) );
 a51533a <=( a51532a  and  a51529a );
 a51534a <=( a51533a  and  a51526a );
 a51537a <=( (not A169)  and  (not A170) );
 a51540a <=( A199  and  (not A168) );
 a51541a <=( a51540a  and  a51537a );
 a51544a <=( A203  and  (not A200) );
 a51547a <=( A233  and  A232 );
 a51548a <=( a51547a  and  a51544a );
 a51549a <=( a51548a  and  a51541a );
 a51552a <=( (not A235)  and  (not A234) );
 a51555a <=( (not A268)  and  (not A267) );
 a51556a <=( a51555a  and  a51552a );
 a51559a <=( (not A298)  and  (not A269) );
 a51562a <=( (not A301)  and  (not A299) );
 a51563a <=( a51562a  and  a51559a );
 a51564a <=( a51563a  and  a51556a );
 a51567a <=( (not A169)  and  (not A170) );
 a51570a <=( A199  and  (not A168) );
 a51571a <=( a51570a  and  a51567a );
 a51574a <=( A203  and  (not A200) );
 a51577a <=( A233  and  A232 );
 a51578a <=( a51577a  and  a51574a );
 a51579a <=( a51578a  and  a51571a );
 a51582a <=( (not A235)  and  (not A234) );
 a51585a <=( (not A266)  and  (not A265) );
 a51586a <=( a51585a  and  a51582a );
 a51589a <=( (not A300)  and  (not A268) );
 a51592a <=( (not A302)  and  (not A301) );
 a51593a <=( a51592a  and  a51589a );
 a51594a <=( a51593a  and  a51586a );
 a51597a <=( (not A169)  and  (not A170) );
 a51600a <=( A199  and  (not A168) );
 a51601a <=( a51600a  and  a51597a );
 a51604a <=( A203  and  (not A200) );
 a51607a <=( A233  and  A232 );
 a51608a <=( a51607a  and  a51604a );
 a51609a <=( a51608a  and  a51601a );
 a51612a <=( (not A235)  and  (not A234) );
 a51615a <=( (not A266)  and  (not A265) );
 a51616a <=( a51615a  and  a51612a );
 a51619a <=( (not A298)  and  (not A268) );
 a51622a <=( (not A301)  and  (not A299) );
 a51623a <=( a51622a  and  a51619a );
 a51624a <=( a51623a  and  a51616a );
 a51627a <=( (not A169)  and  (not A170) );
 a51630a <=( A199  and  (not A168) );
 a51631a <=( a51630a  and  a51627a );
 a51634a <=( A203  and  (not A200) );
 a51637a <=( (not A233)  and  (not A232) );
 a51638a <=( a51637a  and  a51634a );
 a51639a <=( a51638a  and  a51631a );
 a51642a <=( (not A267)  and  (not A235) );
 a51645a <=( (not A269)  and  (not A268) );
 a51646a <=( a51645a  and  a51642a );
 a51649a <=( A299  and  A298 );
 a51652a <=( (not A301)  and  (not A300) );
 a51653a <=( a51652a  and  a51649a );
 a51654a <=( a51653a  and  a51646a );
 a51657a <=( (not A169)  and  (not A170) );
 a51660a <=( A199  and  (not A168) );
 a51661a <=( a51660a  and  a51657a );
 a51664a <=( A203  and  (not A200) );
 a51667a <=( (not A233)  and  (not A232) );
 a51668a <=( a51667a  and  a51664a );
 a51669a <=( a51668a  and  a51661a );
 a51672a <=( A265  and  (not A235) );
 a51675a <=( (not A267)  and  A266 );
 a51676a <=( a51675a  and  a51672a );
 a51679a <=( (not A300)  and  (not A268) );
 a51682a <=( (not A302)  and  (not A301) );
 a51683a <=( a51682a  and  a51679a );
 a51684a <=( a51683a  and  a51676a );
 a51687a <=( (not A169)  and  (not A170) );
 a51690a <=( A199  and  (not A168) );
 a51691a <=( a51690a  and  a51687a );
 a51694a <=( A203  and  (not A200) );
 a51697a <=( (not A233)  and  (not A232) );
 a51698a <=( a51697a  and  a51694a );
 a51699a <=( a51698a  and  a51691a );
 a51702a <=( A265  and  (not A235) );
 a51705a <=( (not A267)  and  A266 );
 a51706a <=( a51705a  and  a51702a );
 a51709a <=( (not A298)  and  (not A268) );
 a51712a <=( (not A301)  and  (not A299) );
 a51713a <=( a51712a  and  a51709a );
 a51714a <=( a51713a  and  a51706a );
 a51717a <=( (not A169)  and  (not A170) );
 a51720a <=( A199  and  (not A168) );
 a51721a <=( a51720a  and  a51717a );
 a51724a <=( A203  and  (not A200) );
 a51727a <=( (not A233)  and  (not A232) );
 a51728a <=( a51727a  and  a51724a );
 a51729a <=( a51728a  and  a51721a );
 a51732a <=( (not A265)  and  (not A235) );
 a51735a <=( (not A268)  and  (not A266) );
 a51736a <=( a51735a  and  a51732a );
 a51739a <=( A299  and  A298 );
 a51742a <=( (not A301)  and  (not A300) );
 a51743a <=( a51742a  and  a51739a );
 a51744a <=( a51743a  and  a51736a );
 a51747a <=( A166  and  A168 );
 a51750a <=( (not A202)  and  (not A201) );
 a51751a <=( a51750a  and  a51747a );
 a51754a <=( A232  and  (not A203) );
 a51757a <=( (not A234)  and  A233 );
 a51758a <=( a51757a  and  a51754a );
 a51759a <=( a51758a  and  a51751a );
 a51762a <=( A265  and  (not A235) );
 a51765a <=( (not A267)  and  A266 );
 a51766a <=( a51765a  and  a51762a );
 a51769a <=( A298  and  (not A268) );
 a51773a <=( (not A301)  and  (not A300) );
 a51774a <=( A299  and  a51773a );
 a51775a <=( a51774a  and  a51769a );
 a51776a <=( a51775a  and  a51766a );
 a51779a <=( A166  and  A168 );
 a51782a <=( A200  and  A199 );
 a51783a <=( a51782a  and  a51779a );
 a51786a <=( (not A202)  and  (not A201) );
 a51789a <=( (not A235)  and  (not A234) );
 a51790a <=( a51789a  and  a51786a );
 a51791a <=( a51790a  and  a51783a );
 a51794a <=( A265  and  (not A236) );
 a51797a <=( (not A267)  and  A266 );
 a51798a <=( a51797a  and  a51794a );
 a51801a <=( A298  and  (not A268) );
 a51805a <=( (not A301)  and  (not A300) );
 a51806a <=( A299  and  a51805a );
 a51807a <=( a51806a  and  a51801a );
 a51808a <=( a51807a  and  a51798a );
 a51811a <=( A166  and  A168 );
 a51814a <=( A200  and  A199 );
 a51815a <=( a51814a  and  a51811a );
 a51818a <=( (not A202)  and  (not A201) );
 a51821a <=( A233  and  A232 );
 a51822a <=( a51821a  and  a51818a );
 a51823a <=( a51822a  and  a51815a );
 a51826a <=( (not A235)  and  (not A234) );
 a51829a <=( (not A268)  and  (not A267) );
 a51830a <=( a51829a  and  a51826a );
 a51833a <=( A298  and  (not A269) );
 a51837a <=( (not A301)  and  (not A300) );
 a51838a <=( A299  and  a51837a );
 a51839a <=( a51838a  and  a51833a );
 a51840a <=( a51839a  and  a51830a );
 a51843a <=( A166  and  A168 );
 a51846a <=( A200  and  A199 );
 a51847a <=( a51846a  and  a51843a );
 a51850a <=( (not A202)  and  (not A201) );
 a51853a <=( A233  and  A232 );
 a51854a <=( a51853a  and  a51850a );
 a51855a <=( a51854a  and  a51847a );
 a51858a <=( (not A235)  and  (not A234) );
 a51861a <=( A266  and  A265 );
 a51862a <=( a51861a  and  a51858a );
 a51865a <=( (not A268)  and  (not A267) );
 a51869a <=( (not A302)  and  (not A301) );
 a51870a <=( (not A300)  and  a51869a );
 a51871a <=( a51870a  and  a51865a );
 a51872a <=( a51871a  and  a51862a );
 a51875a <=( A166  and  A168 );
 a51878a <=( A200  and  A199 );
 a51879a <=( a51878a  and  a51875a );
 a51882a <=( (not A202)  and  (not A201) );
 a51885a <=( A233  and  A232 );
 a51886a <=( a51885a  and  a51882a );
 a51887a <=( a51886a  and  a51879a );
 a51890a <=( (not A235)  and  (not A234) );
 a51893a <=( A266  and  A265 );
 a51894a <=( a51893a  and  a51890a );
 a51897a <=( (not A268)  and  (not A267) );
 a51901a <=( (not A301)  and  (not A299) );
 a51902a <=( (not A298)  and  a51901a );
 a51903a <=( a51902a  and  a51897a );
 a51904a <=( a51903a  and  a51894a );
 a51907a <=( A166  and  A168 );
 a51910a <=( A200  and  A199 );
 a51911a <=( a51910a  and  a51907a );
 a51914a <=( (not A202)  and  (not A201) );
 a51917a <=( A233  and  A232 );
 a51918a <=( a51917a  and  a51914a );
 a51919a <=( a51918a  and  a51911a );
 a51922a <=( (not A235)  and  (not A234) );
 a51925a <=( (not A266)  and  (not A265) );
 a51926a <=( a51925a  and  a51922a );
 a51929a <=( A298  and  (not A268) );
 a51933a <=( (not A301)  and  (not A300) );
 a51934a <=( A299  and  a51933a );
 a51935a <=( a51934a  and  a51929a );
 a51936a <=( a51935a  and  a51926a );
 a51939a <=( A166  and  A168 );
 a51942a <=( A200  and  A199 );
 a51943a <=( a51942a  and  a51939a );
 a51946a <=( (not A202)  and  (not A201) );
 a51949a <=( (not A233)  and  (not A232) );
 a51950a <=( a51949a  and  a51946a );
 a51951a <=( a51950a  and  a51943a );
 a51954a <=( A265  and  (not A235) );
 a51957a <=( (not A267)  and  A266 );
 a51958a <=( a51957a  and  a51954a );
 a51961a <=( A298  and  (not A268) );
 a51965a <=( (not A301)  and  (not A300) );
 a51966a <=( A299  and  a51965a );
 a51967a <=( a51966a  and  a51961a );
 a51968a <=( a51967a  and  a51958a );
 a51971a <=( A166  and  A168 );
 a51974a <=( (not A200)  and  (not A199) );
 a51975a <=( a51974a  and  a51971a );
 a51978a <=( A232  and  (not A202) );
 a51981a <=( (not A234)  and  A233 );
 a51982a <=( a51981a  and  a51978a );
 a51983a <=( a51982a  and  a51975a );
 a51986a <=( A265  and  (not A235) );
 a51989a <=( (not A267)  and  A266 );
 a51990a <=( a51989a  and  a51986a );
 a51993a <=( A298  and  (not A268) );
 a51997a <=( (not A301)  and  (not A300) );
 a51998a <=( A299  and  a51997a );
 a51999a <=( a51998a  and  a51993a );
 a52000a <=( a51999a  and  a51990a );
 a52003a <=( A167  and  A168 );
 a52006a <=( (not A202)  and  (not A201) );
 a52007a <=( a52006a  and  a52003a );
 a52010a <=( A232  and  (not A203) );
 a52013a <=( (not A234)  and  A233 );
 a52014a <=( a52013a  and  a52010a );
 a52015a <=( a52014a  and  a52007a );
 a52018a <=( A265  and  (not A235) );
 a52021a <=( (not A267)  and  A266 );
 a52022a <=( a52021a  and  a52018a );
 a52025a <=( A298  and  (not A268) );
 a52029a <=( (not A301)  and  (not A300) );
 a52030a <=( A299  and  a52029a );
 a52031a <=( a52030a  and  a52025a );
 a52032a <=( a52031a  and  a52022a );
 a52035a <=( A167  and  A168 );
 a52038a <=( A200  and  A199 );
 a52039a <=( a52038a  and  a52035a );
 a52042a <=( (not A202)  and  (not A201) );
 a52045a <=( (not A235)  and  (not A234) );
 a52046a <=( a52045a  and  a52042a );
 a52047a <=( a52046a  and  a52039a );
 a52050a <=( A265  and  (not A236) );
 a52053a <=( (not A267)  and  A266 );
 a52054a <=( a52053a  and  a52050a );
 a52057a <=( A298  and  (not A268) );
 a52061a <=( (not A301)  and  (not A300) );
 a52062a <=( A299  and  a52061a );
 a52063a <=( a52062a  and  a52057a );
 a52064a <=( a52063a  and  a52054a );
 a52067a <=( A167  and  A168 );
 a52070a <=( A200  and  A199 );
 a52071a <=( a52070a  and  a52067a );
 a52074a <=( (not A202)  and  (not A201) );
 a52077a <=( A233  and  A232 );
 a52078a <=( a52077a  and  a52074a );
 a52079a <=( a52078a  and  a52071a );
 a52082a <=( (not A235)  and  (not A234) );
 a52085a <=( (not A268)  and  (not A267) );
 a52086a <=( a52085a  and  a52082a );
 a52089a <=( A298  and  (not A269) );
 a52093a <=( (not A301)  and  (not A300) );
 a52094a <=( A299  and  a52093a );
 a52095a <=( a52094a  and  a52089a );
 a52096a <=( a52095a  and  a52086a );
 a52099a <=( A167  and  A168 );
 a52102a <=( A200  and  A199 );
 a52103a <=( a52102a  and  a52099a );
 a52106a <=( (not A202)  and  (not A201) );
 a52109a <=( A233  and  A232 );
 a52110a <=( a52109a  and  a52106a );
 a52111a <=( a52110a  and  a52103a );
 a52114a <=( (not A235)  and  (not A234) );
 a52117a <=( A266  and  A265 );
 a52118a <=( a52117a  and  a52114a );
 a52121a <=( (not A268)  and  (not A267) );
 a52125a <=( (not A302)  and  (not A301) );
 a52126a <=( (not A300)  and  a52125a );
 a52127a <=( a52126a  and  a52121a );
 a52128a <=( a52127a  and  a52118a );
 a52131a <=( A167  and  A168 );
 a52134a <=( A200  and  A199 );
 a52135a <=( a52134a  and  a52131a );
 a52138a <=( (not A202)  and  (not A201) );
 a52141a <=( A233  and  A232 );
 a52142a <=( a52141a  and  a52138a );
 a52143a <=( a52142a  and  a52135a );
 a52146a <=( (not A235)  and  (not A234) );
 a52149a <=( A266  and  A265 );
 a52150a <=( a52149a  and  a52146a );
 a52153a <=( (not A268)  and  (not A267) );
 a52157a <=( (not A301)  and  (not A299) );
 a52158a <=( (not A298)  and  a52157a );
 a52159a <=( a52158a  and  a52153a );
 a52160a <=( a52159a  and  a52150a );
 a52163a <=( A167  and  A168 );
 a52166a <=( A200  and  A199 );
 a52167a <=( a52166a  and  a52163a );
 a52170a <=( (not A202)  and  (not A201) );
 a52173a <=( A233  and  A232 );
 a52174a <=( a52173a  and  a52170a );
 a52175a <=( a52174a  and  a52167a );
 a52178a <=( (not A235)  and  (not A234) );
 a52181a <=( (not A266)  and  (not A265) );
 a52182a <=( a52181a  and  a52178a );
 a52185a <=( A298  and  (not A268) );
 a52189a <=( (not A301)  and  (not A300) );
 a52190a <=( A299  and  a52189a );
 a52191a <=( a52190a  and  a52185a );
 a52192a <=( a52191a  and  a52182a );
 a52195a <=( A167  and  A168 );
 a52198a <=( A200  and  A199 );
 a52199a <=( a52198a  and  a52195a );
 a52202a <=( (not A202)  and  (not A201) );
 a52205a <=( (not A233)  and  (not A232) );
 a52206a <=( a52205a  and  a52202a );
 a52207a <=( a52206a  and  a52199a );
 a52210a <=( A265  and  (not A235) );
 a52213a <=( (not A267)  and  A266 );
 a52214a <=( a52213a  and  a52210a );
 a52217a <=( A298  and  (not A268) );
 a52221a <=( (not A301)  and  (not A300) );
 a52222a <=( A299  and  a52221a );
 a52223a <=( a52222a  and  a52217a );
 a52224a <=( a52223a  and  a52214a );
 a52227a <=( A167  and  A168 );
 a52230a <=( (not A200)  and  (not A199) );
 a52231a <=( a52230a  and  a52227a );
 a52234a <=( A232  and  (not A202) );
 a52237a <=( (not A234)  and  A233 );
 a52238a <=( a52237a  and  a52234a );
 a52239a <=( a52238a  and  a52231a );
 a52242a <=( A265  and  (not A235) );
 a52245a <=( (not A267)  and  A266 );
 a52246a <=( a52245a  and  a52242a );
 a52249a <=( A298  and  (not A268) );
 a52253a <=( (not A301)  and  (not A300) );
 a52254a <=( A299  and  a52253a );
 a52255a <=( a52254a  and  a52249a );
 a52256a <=( a52255a  and  a52246a );
 a52259a <=( A167  and  A170 );
 a52262a <=( (not A201)  and  (not A166) );
 a52263a <=( a52262a  and  a52259a );
 a52266a <=( (not A203)  and  (not A202) );
 a52269a <=( (not A235)  and  (not A234) );
 a52270a <=( a52269a  and  a52266a );
 a52271a <=( a52270a  and  a52263a );
 a52274a <=( A265  and  (not A236) );
 a52277a <=( (not A267)  and  A266 );
 a52278a <=( a52277a  and  a52274a );
 a52281a <=( A298  and  (not A268) );
 a52285a <=( (not A301)  and  (not A300) );
 a52286a <=( A299  and  a52285a );
 a52287a <=( a52286a  and  a52281a );
 a52288a <=( a52287a  and  a52278a );
 a52291a <=( A167  and  A170 );
 a52294a <=( (not A201)  and  (not A166) );
 a52295a <=( a52294a  and  a52291a );
 a52298a <=( (not A203)  and  (not A202) );
 a52301a <=( A233  and  A232 );
 a52302a <=( a52301a  and  a52298a );
 a52303a <=( a52302a  and  a52295a );
 a52306a <=( (not A235)  and  (not A234) );
 a52309a <=( (not A268)  and  (not A267) );
 a52310a <=( a52309a  and  a52306a );
 a52313a <=( A298  and  (not A269) );
 a52317a <=( (not A301)  and  (not A300) );
 a52318a <=( A299  and  a52317a );
 a52319a <=( a52318a  and  a52313a );
 a52320a <=( a52319a  and  a52310a );
 a52323a <=( A167  and  A170 );
 a52326a <=( (not A201)  and  (not A166) );
 a52327a <=( a52326a  and  a52323a );
 a52330a <=( (not A203)  and  (not A202) );
 a52333a <=( A233  and  A232 );
 a52334a <=( a52333a  and  a52330a );
 a52335a <=( a52334a  and  a52327a );
 a52338a <=( (not A235)  and  (not A234) );
 a52341a <=( A266  and  A265 );
 a52342a <=( a52341a  and  a52338a );
 a52345a <=( (not A268)  and  (not A267) );
 a52349a <=( (not A302)  and  (not A301) );
 a52350a <=( (not A300)  and  a52349a );
 a52351a <=( a52350a  and  a52345a );
 a52352a <=( a52351a  and  a52342a );
 a52355a <=( A167  and  A170 );
 a52358a <=( (not A201)  and  (not A166) );
 a52359a <=( a52358a  and  a52355a );
 a52362a <=( (not A203)  and  (not A202) );
 a52365a <=( A233  and  A232 );
 a52366a <=( a52365a  and  a52362a );
 a52367a <=( a52366a  and  a52359a );
 a52370a <=( (not A235)  and  (not A234) );
 a52373a <=( A266  and  A265 );
 a52374a <=( a52373a  and  a52370a );
 a52377a <=( (not A268)  and  (not A267) );
 a52381a <=( (not A301)  and  (not A299) );
 a52382a <=( (not A298)  and  a52381a );
 a52383a <=( a52382a  and  a52377a );
 a52384a <=( a52383a  and  a52374a );
 a52387a <=( A167  and  A170 );
 a52390a <=( (not A201)  and  (not A166) );
 a52391a <=( a52390a  and  a52387a );
 a52394a <=( (not A203)  and  (not A202) );
 a52397a <=( A233  and  A232 );
 a52398a <=( a52397a  and  a52394a );
 a52399a <=( a52398a  and  a52391a );
 a52402a <=( (not A235)  and  (not A234) );
 a52405a <=( (not A266)  and  (not A265) );
 a52406a <=( a52405a  and  a52402a );
 a52409a <=( A298  and  (not A268) );
 a52413a <=( (not A301)  and  (not A300) );
 a52414a <=( A299  and  a52413a );
 a52415a <=( a52414a  and  a52409a );
 a52416a <=( a52415a  and  a52406a );
 a52419a <=( A167  and  A170 );
 a52422a <=( (not A201)  and  (not A166) );
 a52423a <=( a52422a  and  a52419a );
 a52426a <=( (not A203)  and  (not A202) );
 a52429a <=( (not A233)  and  (not A232) );
 a52430a <=( a52429a  and  a52426a );
 a52431a <=( a52430a  and  a52423a );
 a52434a <=( A265  and  (not A235) );
 a52437a <=( (not A267)  and  A266 );
 a52438a <=( a52437a  and  a52434a );
 a52441a <=( A298  and  (not A268) );
 a52445a <=( (not A301)  and  (not A300) );
 a52446a <=( A299  and  a52445a );
 a52447a <=( a52446a  and  a52441a );
 a52448a <=( a52447a  and  a52438a );
 a52451a <=( A167  and  A170 );
 a52454a <=( A199  and  (not A166) );
 a52455a <=( a52454a  and  a52451a );
 a52458a <=( (not A201)  and  A200 );
 a52461a <=( (not A234)  and  (not A202) );
 a52462a <=( a52461a  and  a52458a );
 a52463a <=( a52462a  and  a52455a );
 a52466a <=( (not A236)  and  (not A235) );
 a52469a <=( (not A268)  and  (not A267) );
 a52470a <=( a52469a  and  a52466a );
 a52473a <=( A298  and  (not A269) );
 a52477a <=( (not A301)  and  (not A300) );
 a52478a <=( A299  and  a52477a );
 a52479a <=( a52478a  and  a52473a );
 a52480a <=( a52479a  and  a52470a );
 a52483a <=( A167  and  A170 );
 a52486a <=( A199  and  (not A166) );
 a52487a <=( a52486a  and  a52483a );
 a52490a <=( (not A201)  and  A200 );
 a52493a <=( (not A234)  and  (not A202) );
 a52494a <=( a52493a  and  a52490a );
 a52495a <=( a52494a  and  a52487a );
 a52498a <=( (not A236)  and  (not A235) );
 a52501a <=( A266  and  A265 );
 a52502a <=( a52501a  and  a52498a );
 a52505a <=( (not A268)  and  (not A267) );
 a52509a <=( (not A302)  and  (not A301) );
 a52510a <=( (not A300)  and  a52509a );
 a52511a <=( a52510a  and  a52505a );
 a52512a <=( a52511a  and  a52502a );
 a52515a <=( A167  and  A170 );
 a52518a <=( A199  and  (not A166) );
 a52519a <=( a52518a  and  a52515a );
 a52522a <=( (not A201)  and  A200 );
 a52525a <=( (not A234)  and  (not A202) );
 a52526a <=( a52525a  and  a52522a );
 a52527a <=( a52526a  and  a52519a );
 a52530a <=( (not A236)  and  (not A235) );
 a52533a <=( A266  and  A265 );
 a52534a <=( a52533a  and  a52530a );
 a52537a <=( (not A268)  and  (not A267) );
 a52541a <=( (not A301)  and  (not A299) );
 a52542a <=( (not A298)  and  a52541a );
 a52543a <=( a52542a  and  a52537a );
 a52544a <=( a52543a  and  a52534a );
 a52547a <=( A167  and  A170 );
 a52550a <=( A199  and  (not A166) );
 a52551a <=( a52550a  and  a52547a );
 a52554a <=( (not A201)  and  A200 );
 a52557a <=( (not A234)  and  (not A202) );
 a52558a <=( a52557a  and  a52554a );
 a52559a <=( a52558a  and  a52551a );
 a52562a <=( (not A236)  and  (not A235) );
 a52565a <=( (not A266)  and  (not A265) );
 a52566a <=( a52565a  and  a52562a );
 a52569a <=( A298  and  (not A268) );
 a52573a <=( (not A301)  and  (not A300) );
 a52574a <=( A299  and  a52573a );
 a52575a <=( a52574a  and  a52569a );
 a52576a <=( a52575a  and  a52566a );
 a52579a <=( A167  and  A170 );
 a52582a <=( A199  and  (not A166) );
 a52583a <=( a52582a  and  a52579a );
 a52586a <=( (not A201)  and  A200 );
 a52589a <=( A232  and  (not A202) );
 a52590a <=( a52589a  and  a52586a );
 a52591a <=( a52590a  and  a52583a );
 a52594a <=( (not A234)  and  A233 );
 a52597a <=( (not A267)  and  (not A235) );
 a52598a <=( a52597a  and  a52594a );
 a52601a <=( (not A269)  and  (not A268) );
 a52605a <=( (not A302)  and  (not A301) );
 a52606a <=( (not A300)  and  a52605a );
 a52607a <=( a52606a  and  a52601a );
 a52608a <=( a52607a  and  a52598a );
 a52611a <=( A167  and  A170 );
 a52614a <=( A199  and  (not A166) );
 a52615a <=( a52614a  and  a52611a );
 a52618a <=( (not A201)  and  A200 );
 a52621a <=( A232  and  (not A202) );
 a52622a <=( a52621a  and  a52618a );
 a52623a <=( a52622a  and  a52615a );
 a52626a <=( (not A234)  and  A233 );
 a52629a <=( (not A267)  and  (not A235) );
 a52630a <=( a52629a  and  a52626a );
 a52633a <=( (not A269)  and  (not A268) );
 a52637a <=( (not A301)  and  (not A299) );
 a52638a <=( (not A298)  and  a52637a );
 a52639a <=( a52638a  and  a52633a );
 a52640a <=( a52639a  and  a52630a );
 a52643a <=( A167  and  A170 );
 a52646a <=( A199  and  (not A166) );
 a52647a <=( a52646a  and  a52643a );
 a52650a <=( (not A201)  and  A200 );
 a52653a <=( A232  and  (not A202) );
 a52654a <=( a52653a  and  a52650a );
 a52655a <=( a52654a  and  a52647a );
 a52658a <=( (not A234)  and  A233 );
 a52661a <=( (not A265)  and  (not A235) );
 a52662a <=( a52661a  and  a52658a );
 a52665a <=( (not A268)  and  (not A266) );
 a52669a <=( (not A302)  and  (not A301) );
 a52670a <=( (not A300)  and  a52669a );
 a52671a <=( a52670a  and  a52665a );
 a52672a <=( a52671a  and  a52662a );
 a52675a <=( A167  and  A170 );
 a52678a <=( A199  and  (not A166) );
 a52679a <=( a52678a  and  a52675a );
 a52682a <=( (not A201)  and  A200 );
 a52685a <=( A232  and  (not A202) );
 a52686a <=( a52685a  and  a52682a );
 a52687a <=( a52686a  and  a52679a );
 a52690a <=( (not A234)  and  A233 );
 a52693a <=( (not A265)  and  (not A235) );
 a52694a <=( a52693a  and  a52690a );
 a52697a <=( (not A268)  and  (not A266) );
 a52701a <=( (not A301)  and  (not A299) );
 a52702a <=( (not A298)  and  a52701a );
 a52703a <=( a52702a  and  a52697a );
 a52704a <=( a52703a  and  a52694a );
 a52707a <=( A167  and  A170 );
 a52710a <=( A199  and  (not A166) );
 a52711a <=( a52710a  and  a52707a );
 a52714a <=( (not A201)  and  A200 );
 a52717a <=( (not A232)  and  (not A202) );
 a52718a <=( a52717a  and  a52714a );
 a52719a <=( a52718a  and  a52711a );
 a52722a <=( (not A235)  and  (not A233) );
 a52725a <=( (not A268)  and  (not A267) );
 a52726a <=( a52725a  and  a52722a );
 a52729a <=( A298  and  (not A269) );
 a52733a <=( (not A301)  and  (not A300) );
 a52734a <=( A299  and  a52733a );
 a52735a <=( a52734a  and  a52729a );
 a52736a <=( a52735a  and  a52726a );
 a52739a <=( A167  and  A170 );
 a52742a <=( A199  and  (not A166) );
 a52743a <=( a52742a  and  a52739a );
 a52746a <=( (not A201)  and  A200 );
 a52749a <=( (not A232)  and  (not A202) );
 a52750a <=( a52749a  and  a52746a );
 a52751a <=( a52750a  and  a52743a );
 a52754a <=( (not A235)  and  (not A233) );
 a52757a <=( A266  and  A265 );
 a52758a <=( a52757a  and  a52754a );
 a52761a <=( (not A268)  and  (not A267) );
 a52765a <=( (not A302)  and  (not A301) );
 a52766a <=( (not A300)  and  a52765a );
 a52767a <=( a52766a  and  a52761a );
 a52768a <=( a52767a  and  a52758a );
 a52771a <=( A167  and  A170 );
 a52774a <=( A199  and  (not A166) );
 a52775a <=( a52774a  and  a52771a );
 a52778a <=( (not A201)  and  A200 );
 a52781a <=( (not A232)  and  (not A202) );
 a52782a <=( a52781a  and  a52778a );
 a52783a <=( a52782a  and  a52775a );
 a52786a <=( (not A235)  and  (not A233) );
 a52789a <=( A266  and  A265 );
 a52790a <=( a52789a  and  a52786a );
 a52793a <=( (not A268)  and  (not A267) );
 a52797a <=( (not A301)  and  (not A299) );
 a52798a <=( (not A298)  and  a52797a );
 a52799a <=( a52798a  and  a52793a );
 a52800a <=( a52799a  and  a52790a );
 a52803a <=( A167  and  A170 );
 a52806a <=( A199  and  (not A166) );
 a52807a <=( a52806a  and  a52803a );
 a52810a <=( (not A201)  and  A200 );
 a52813a <=( (not A232)  and  (not A202) );
 a52814a <=( a52813a  and  a52810a );
 a52815a <=( a52814a  and  a52807a );
 a52818a <=( (not A235)  and  (not A233) );
 a52821a <=( (not A266)  and  (not A265) );
 a52822a <=( a52821a  and  a52818a );
 a52825a <=( A298  and  (not A268) );
 a52829a <=( (not A301)  and  (not A300) );
 a52830a <=( A299  and  a52829a );
 a52831a <=( a52830a  and  a52825a );
 a52832a <=( a52831a  and  a52822a );
 a52835a <=( A167  and  A170 );
 a52838a <=( (not A199)  and  (not A166) );
 a52839a <=( a52838a  and  a52835a );
 a52842a <=( (not A202)  and  (not A200) );
 a52845a <=( (not A235)  and  (not A234) );
 a52846a <=( a52845a  and  a52842a );
 a52847a <=( a52846a  and  a52839a );
 a52850a <=( A265  and  (not A236) );
 a52853a <=( (not A267)  and  A266 );
 a52854a <=( a52853a  and  a52850a );
 a52857a <=( A298  and  (not A268) );
 a52861a <=( (not A301)  and  (not A300) );
 a52862a <=( A299  and  a52861a );
 a52863a <=( a52862a  and  a52857a );
 a52864a <=( a52863a  and  a52854a );
 a52867a <=( A167  and  A170 );
 a52870a <=( (not A199)  and  (not A166) );
 a52871a <=( a52870a  and  a52867a );
 a52874a <=( (not A202)  and  (not A200) );
 a52877a <=( A233  and  A232 );
 a52878a <=( a52877a  and  a52874a );
 a52879a <=( a52878a  and  a52871a );
 a52882a <=( (not A235)  and  (not A234) );
 a52885a <=( (not A268)  and  (not A267) );
 a52886a <=( a52885a  and  a52882a );
 a52889a <=( A298  and  (not A269) );
 a52893a <=( (not A301)  and  (not A300) );
 a52894a <=( A299  and  a52893a );
 a52895a <=( a52894a  and  a52889a );
 a52896a <=( a52895a  and  a52886a );
 a52899a <=( A167  and  A170 );
 a52902a <=( (not A199)  and  (not A166) );
 a52903a <=( a52902a  and  a52899a );
 a52906a <=( (not A202)  and  (not A200) );
 a52909a <=( A233  and  A232 );
 a52910a <=( a52909a  and  a52906a );
 a52911a <=( a52910a  and  a52903a );
 a52914a <=( (not A235)  and  (not A234) );
 a52917a <=( A266  and  A265 );
 a52918a <=( a52917a  and  a52914a );
 a52921a <=( (not A268)  and  (not A267) );
 a52925a <=( (not A302)  and  (not A301) );
 a52926a <=( (not A300)  and  a52925a );
 a52927a <=( a52926a  and  a52921a );
 a52928a <=( a52927a  and  a52918a );
 a52931a <=( A167  and  A170 );
 a52934a <=( (not A199)  and  (not A166) );
 a52935a <=( a52934a  and  a52931a );
 a52938a <=( (not A202)  and  (not A200) );
 a52941a <=( A233  and  A232 );
 a52942a <=( a52941a  and  a52938a );
 a52943a <=( a52942a  and  a52935a );
 a52946a <=( (not A235)  and  (not A234) );
 a52949a <=( A266  and  A265 );
 a52950a <=( a52949a  and  a52946a );
 a52953a <=( (not A268)  and  (not A267) );
 a52957a <=( (not A301)  and  (not A299) );
 a52958a <=( (not A298)  and  a52957a );
 a52959a <=( a52958a  and  a52953a );
 a52960a <=( a52959a  and  a52950a );
 a52963a <=( A167  and  A170 );
 a52966a <=( (not A199)  and  (not A166) );
 a52967a <=( a52966a  and  a52963a );
 a52970a <=( (not A202)  and  (not A200) );
 a52973a <=( A233  and  A232 );
 a52974a <=( a52973a  and  a52970a );
 a52975a <=( a52974a  and  a52967a );
 a52978a <=( (not A235)  and  (not A234) );
 a52981a <=( (not A266)  and  (not A265) );
 a52982a <=( a52981a  and  a52978a );
 a52985a <=( A298  and  (not A268) );
 a52989a <=( (not A301)  and  (not A300) );
 a52990a <=( A299  and  a52989a );
 a52991a <=( a52990a  and  a52985a );
 a52992a <=( a52991a  and  a52982a );
 a52995a <=( A167  and  A170 );
 a52998a <=( (not A199)  and  (not A166) );
 a52999a <=( a52998a  and  a52995a );
 a53002a <=( (not A202)  and  (not A200) );
 a53005a <=( (not A233)  and  (not A232) );
 a53006a <=( a53005a  and  a53002a );
 a53007a <=( a53006a  and  a52999a );
 a53010a <=( A265  and  (not A235) );
 a53013a <=( (not A267)  and  A266 );
 a53014a <=( a53013a  and  a53010a );
 a53017a <=( A298  and  (not A268) );
 a53021a <=( (not A301)  and  (not A300) );
 a53022a <=( A299  and  a53021a );
 a53023a <=( a53022a  and  a53017a );
 a53024a <=( a53023a  and  a53014a );
 a53027a <=( (not A167)  and  A170 );
 a53030a <=( (not A201)  and  A166 );
 a53031a <=( a53030a  and  a53027a );
 a53034a <=( (not A203)  and  (not A202) );
 a53037a <=( (not A235)  and  (not A234) );
 a53038a <=( a53037a  and  a53034a );
 a53039a <=( a53038a  and  a53031a );
 a53042a <=( A265  and  (not A236) );
 a53045a <=( (not A267)  and  A266 );
 a53046a <=( a53045a  and  a53042a );
 a53049a <=( A298  and  (not A268) );
 a53053a <=( (not A301)  and  (not A300) );
 a53054a <=( A299  and  a53053a );
 a53055a <=( a53054a  and  a53049a );
 a53056a <=( a53055a  and  a53046a );
 a53059a <=( (not A167)  and  A170 );
 a53062a <=( (not A201)  and  A166 );
 a53063a <=( a53062a  and  a53059a );
 a53066a <=( (not A203)  and  (not A202) );
 a53069a <=( A233  and  A232 );
 a53070a <=( a53069a  and  a53066a );
 a53071a <=( a53070a  and  a53063a );
 a53074a <=( (not A235)  and  (not A234) );
 a53077a <=( (not A268)  and  (not A267) );
 a53078a <=( a53077a  and  a53074a );
 a53081a <=( A298  and  (not A269) );
 a53085a <=( (not A301)  and  (not A300) );
 a53086a <=( A299  and  a53085a );
 a53087a <=( a53086a  and  a53081a );
 a53088a <=( a53087a  and  a53078a );
 a53091a <=( (not A167)  and  A170 );
 a53094a <=( (not A201)  and  A166 );
 a53095a <=( a53094a  and  a53091a );
 a53098a <=( (not A203)  and  (not A202) );
 a53101a <=( A233  and  A232 );
 a53102a <=( a53101a  and  a53098a );
 a53103a <=( a53102a  and  a53095a );
 a53106a <=( (not A235)  and  (not A234) );
 a53109a <=( A266  and  A265 );
 a53110a <=( a53109a  and  a53106a );
 a53113a <=( (not A268)  and  (not A267) );
 a53117a <=( (not A302)  and  (not A301) );
 a53118a <=( (not A300)  and  a53117a );
 a53119a <=( a53118a  and  a53113a );
 a53120a <=( a53119a  and  a53110a );
 a53123a <=( (not A167)  and  A170 );
 a53126a <=( (not A201)  and  A166 );
 a53127a <=( a53126a  and  a53123a );
 a53130a <=( (not A203)  and  (not A202) );
 a53133a <=( A233  and  A232 );
 a53134a <=( a53133a  and  a53130a );
 a53135a <=( a53134a  and  a53127a );
 a53138a <=( (not A235)  and  (not A234) );
 a53141a <=( A266  and  A265 );
 a53142a <=( a53141a  and  a53138a );
 a53145a <=( (not A268)  and  (not A267) );
 a53149a <=( (not A301)  and  (not A299) );
 a53150a <=( (not A298)  and  a53149a );
 a53151a <=( a53150a  and  a53145a );
 a53152a <=( a53151a  and  a53142a );
 a53155a <=( (not A167)  and  A170 );
 a53158a <=( (not A201)  and  A166 );
 a53159a <=( a53158a  and  a53155a );
 a53162a <=( (not A203)  and  (not A202) );
 a53165a <=( A233  and  A232 );
 a53166a <=( a53165a  and  a53162a );
 a53167a <=( a53166a  and  a53159a );
 a53170a <=( (not A235)  and  (not A234) );
 a53173a <=( (not A266)  and  (not A265) );
 a53174a <=( a53173a  and  a53170a );
 a53177a <=( A298  and  (not A268) );
 a53181a <=( (not A301)  and  (not A300) );
 a53182a <=( A299  and  a53181a );
 a53183a <=( a53182a  and  a53177a );
 a53184a <=( a53183a  and  a53174a );
 a53187a <=( (not A167)  and  A170 );
 a53190a <=( (not A201)  and  A166 );
 a53191a <=( a53190a  and  a53187a );
 a53194a <=( (not A203)  and  (not A202) );
 a53197a <=( (not A233)  and  (not A232) );
 a53198a <=( a53197a  and  a53194a );
 a53199a <=( a53198a  and  a53191a );
 a53202a <=( A265  and  (not A235) );
 a53205a <=( (not A267)  and  A266 );
 a53206a <=( a53205a  and  a53202a );
 a53209a <=( A298  and  (not A268) );
 a53213a <=( (not A301)  and  (not A300) );
 a53214a <=( A299  and  a53213a );
 a53215a <=( a53214a  and  a53209a );
 a53216a <=( a53215a  and  a53206a );
 a53219a <=( (not A167)  and  A170 );
 a53222a <=( A199  and  A166 );
 a53223a <=( a53222a  and  a53219a );
 a53226a <=( (not A201)  and  A200 );
 a53229a <=( (not A234)  and  (not A202) );
 a53230a <=( a53229a  and  a53226a );
 a53231a <=( a53230a  and  a53223a );
 a53234a <=( (not A236)  and  (not A235) );
 a53237a <=( (not A268)  and  (not A267) );
 a53238a <=( a53237a  and  a53234a );
 a53241a <=( A298  and  (not A269) );
 a53245a <=( (not A301)  and  (not A300) );
 a53246a <=( A299  and  a53245a );
 a53247a <=( a53246a  and  a53241a );
 a53248a <=( a53247a  and  a53238a );
 a53251a <=( (not A167)  and  A170 );
 a53254a <=( A199  and  A166 );
 a53255a <=( a53254a  and  a53251a );
 a53258a <=( (not A201)  and  A200 );
 a53261a <=( (not A234)  and  (not A202) );
 a53262a <=( a53261a  and  a53258a );
 a53263a <=( a53262a  and  a53255a );
 a53266a <=( (not A236)  and  (not A235) );
 a53269a <=( A266  and  A265 );
 a53270a <=( a53269a  and  a53266a );
 a53273a <=( (not A268)  and  (not A267) );
 a53277a <=( (not A302)  and  (not A301) );
 a53278a <=( (not A300)  and  a53277a );
 a53279a <=( a53278a  and  a53273a );
 a53280a <=( a53279a  and  a53270a );
 a53283a <=( (not A167)  and  A170 );
 a53286a <=( A199  and  A166 );
 a53287a <=( a53286a  and  a53283a );
 a53290a <=( (not A201)  and  A200 );
 a53293a <=( (not A234)  and  (not A202) );
 a53294a <=( a53293a  and  a53290a );
 a53295a <=( a53294a  and  a53287a );
 a53298a <=( (not A236)  and  (not A235) );
 a53301a <=( A266  and  A265 );
 a53302a <=( a53301a  and  a53298a );
 a53305a <=( (not A268)  and  (not A267) );
 a53309a <=( (not A301)  and  (not A299) );
 a53310a <=( (not A298)  and  a53309a );
 a53311a <=( a53310a  and  a53305a );
 a53312a <=( a53311a  and  a53302a );
 a53315a <=( (not A167)  and  A170 );
 a53318a <=( A199  and  A166 );
 a53319a <=( a53318a  and  a53315a );
 a53322a <=( (not A201)  and  A200 );
 a53325a <=( (not A234)  and  (not A202) );
 a53326a <=( a53325a  and  a53322a );
 a53327a <=( a53326a  and  a53319a );
 a53330a <=( (not A236)  and  (not A235) );
 a53333a <=( (not A266)  and  (not A265) );
 a53334a <=( a53333a  and  a53330a );
 a53337a <=( A298  and  (not A268) );
 a53341a <=( (not A301)  and  (not A300) );
 a53342a <=( A299  and  a53341a );
 a53343a <=( a53342a  and  a53337a );
 a53344a <=( a53343a  and  a53334a );
 a53347a <=( (not A167)  and  A170 );
 a53350a <=( A199  and  A166 );
 a53351a <=( a53350a  and  a53347a );
 a53354a <=( (not A201)  and  A200 );
 a53357a <=( A232  and  (not A202) );
 a53358a <=( a53357a  and  a53354a );
 a53359a <=( a53358a  and  a53351a );
 a53362a <=( (not A234)  and  A233 );
 a53365a <=( (not A267)  and  (not A235) );
 a53366a <=( a53365a  and  a53362a );
 a53369a <=( (not A269)  and  (not A268) );
 a53373a <=( (not A302)  and  (not A301) );
 a53374a <=( (not A300)  and  a53373a );
 a53375a <=( a53374a  and  a53369a );
 a53376a <=( a53375a  and  a53366a );
 a53379a <=( (not A167)  and  A170 );
 a53382a <=( A199  and  A166 );
 a53383a <=( a53382a  and  a53379a );
 a53386a <=( (not A201)  and  A200 );
 a53389a <=( A232  and  (not A202) );
 a53390a <=( a53389a  and  a53386a );
 a53391a <=( a53390a  and  a53383a );
 a53394a <=( (not A234)  and  A233 );
 a53397a <=( (not A267)  and  (not A235) );
 a53398a <=( a53397a  and  a53394a );
 a53401a <=( (not A269)  and  (not A268) );
 a53405a <=( (not A301)  and  (not A299) );
 a53406a <=( (not A298)  and  a53405a );
 a53407a <=( a53406a  and  a53401a );
 a53408a <=( a53407a  and  a53398a );
 a53411a <=( (not A167)  and  A170 );
 a53414a <=( A199  and  A166 );
 a53415a <=( a53414a  and  a53411a );
 a53418a <=( (not A201)  and  A200 );
 a53421a <=( A232  and  (not A202) );
 a53422a <=( a53421a  and  a53418a );
 a53423a <=( a53422a  and  a53415a );
 a53426a <=( (not A234)  and  A233 );
 a53429a <=( (not A265)  and  (not A235) );
 a53430a <=( a53429a  and  a53426a );
 a53433a <=( (not A268)  and  (not A266) );
 a53437a <=( (not A302)  and  (not A301) );
 a53438a <=( (not A300)  and  a53437a );
 a53439a <=( a53438a  and  a53433a );
 a53440a <=( a53439a  and  a53430a );
 a53443a <=( (not A167)  and  A170 );
 a53446a <=( A199  and  A166 );
 a53447a <=( a53446a  and  a53443a );
 a53450a <=( (not A201)  and  A200 );
 a53453a <=( A232  and  (not A202) );
 a53454a <=( a53453a  and  a53450a );
 a53455a <=( a53454a  and  a53447a );
 a53458a <=( (not A234)  and  A233 );
 a53461a <=( (not A265)  and  (not A235) );
 a53462a <=( a53461a  and  a53458a );
 a53465a <=( (not A268)  and  (not A266) );
 a53469a <=( (not A301)  and  (not A299) );
 a53470a <=( (not A298)  and  a53469a );
 a53471a <=( a53470a  and  a53465a );
 a53472a <=( a53471a  and  a53462a );
 a53475a <=( (not A167)  and  A170 );
 a53478a <=( A199  and  A166 );
 a53479a <=( a53478a  and  a53475a );
 a53482a <=( (not A201)  and  A200 );
 a53485a <=( (not A232)  and  (not A202) );
 a53486a <=( a53485a  and  a53482a );
 a53487a <=( a53486a  and  a53479a );
 a53490a <=( (not A235)  and  (not A233) );
 a53493a <=( (not A268)  and  (not A267) );
 a53494a <=( a53493a  and  a53490a );
 a53497a <=( A298  and  (not A269) );
 a53501a <=( (not A301)  and  (not A300) );
 a53502a <=( A299  and  a53501a );
 a53503a <=( a53502a  and  a53497a );
 a53504a <=( a53503a  and  a53494a );
 a53507a <=( (not A167)  and  A170 );
 a53510a <=( A199  and  A166 );
 a53511a <=( a53510a  and  a53507a );
 a53514a <=( (not A201)  and  A200 );
 a53517a <=( (not A232)  and  (not A202) );
 a53518a <=( a53517a  and  a53514a );
 a53519a <=( a53518a  and  a53511a );
 a53522a <=( (not A235)  and  (not A233) );
 a53525a <=( A266  and  A265 );
 a53526a <=( a53525a  and  a53522a );
 a53529a <=( (not A268)  and  (not A267) );
 a53533a <=( (not A302)  and  (not A301) );
 a53534a <=( (not A300)  and  a53533a );
 a53535a <=( a53534a  and  a53529a );
 a53536a <=( a53535a  and  a53526a );
 a53539a <=( (not A167)  and  A170 );
 a53542a <=( A199  and  A166 );
 a53543a <=( a53542a  and  a53539a );
 a53546a <=( (not A201)  and  A200 );
 a53549a <=( (not A232)  and  (not A202) );
 a53550a <=( a53549a  and  a53546a );
 a53551a <=( a53550a  and  a53543a );
 a53554a <=( (not A235)  and  (not A233) );
 a53557a <=( A266  and  A265 );
 a53558a <=( a53557a  and  a53554a );
 a53561a <=( (not A268)  and  (not A267) );
 a53565a <=( (not A301)  and  (not A299) );
 a53566a <=( (not A298)  and  a53565a );
 a53567a <=( a53566a  and  a53561a );
 a53568a <=( a53567a  and  a53558a );
 a53571a <=( (not A167)  and  A170 );
 a53574a <=( A199  and  A166 );
 a53575a <=( a53574a  and  a53571a );
 a53578a <=( (not A201)  and  A200 );
 a53581a <=( (not A232)  and  (not A202) );
 a53582a <=( a53581a  and  a53578a );
 a53583a <=( a53582a  and  a53575a );
 a53586a <=( (not A235)  and  (not A233) );
 a53589a <=( (not A266)  and  (not A265) );
 a53590a <=( a53589a  and  a53586a );
 a53593a <=( A298  and  (not A268) );
 a53597a <=( (not A301)  and  (not A300) );
 a53598a <=( A299  and  a53597a );
 a53599a <=( a53598a  and  a53593a );
 a53600a <=( a53599a  and  a53590a );
 a53603a <=( (not A167)  and  A170 );
 a53606a <=( (not A199)  and  A166 );
 a53607a <=( a53606a  and  a53603a );
 a53610a <=( (not A202)  and  (not A200) );
 a53613a <=( (not A235)  and  (not A234) );
 a53614a <=( a53613a  and  a53610a );
 a53615a <=( a53614a  and  a53607a );
 a53618a <=( A265  and  (not A236) );
 a53621a <=( (not A267)  and  A266 );
 a53622a <=( a53621a  and  a53618a );
 a53625a <=( A298  and  (not A268) );
 a53629a <=( (not A301)  and  (not A300) );
 a53630a <=( A299  and  a53629a );
 a53631a <=( a53630a  and  a53625a );
 a53632a <=( a53631a  and  a53622a );
 a53635a <=( (not A167)  and  A170 );
 a53638a <=( (not A199)  and  A166 );
 a53639a <=( a53638a  and  a53635a );
 a53642a <=( (not A202)  and  (not A200) );
 a53645a <=( A233  and  A232 );
 a53646a <=( a53645a  and  a53642a );
 a53647a <=( a53646a  and  a53639a );
 a53650a <=( (not A235)  and  (not A234) );
 a53653a <=( (not A268)  and  (not A267) );
 a53654a <=( a53653a  and  a53650a );
 a53657a <=( A298  and  (not A269) );
 a53661a <=( (not A301)  and  (not A300) );
 a53662a <=( A299  and  a53661a );
 a53663a <=( a53662a  and  a53657a );
 a53664a <=( a53663a  and  a53654a );
 a53667a <=( (not A167)  and  A170 );
 a53670a <=( (not A199)  and  A166 );
 a53671a <=( a53670a  and  a53667a );
 a53674a <=( (not A202)  and  (not A200) );
 a53677a <=( A233  and  A232 );
 a53678a <=( a53677a  and  a53674a );
 a53679a <=( a53678a  and  a53671a );
 a53682a <=( (not A235)  and  (not A234) );
 a53685a <=( A266  and  A265 );
 a53686a <=( a53685a  and  a53682a );
 a53689a <=( (not A268)  and  (not A267) );
 a53693a <=( (not A302)  and  (not A301) );
 a53694a <=( (not A300)  and  a53693a );
 a53695a <=( a53694a  and  a53689a );
 a53696a <=( a53695a  and  a53686a );
 a53699a <=( (not A167)  and  A170 );
 a53702a <=( (not A199)  and  A166 );
 a53703a <=( a53702a  and  a53699a );
 a53706a <=( (not A202)  and  (not A200) );
 a53709a <=( A233  and  A232 );
 a53710a <=( a53709a  and  a53706a );
 a53711a <=( a53710a  and  a53703a );
 a53714a <=( (not A235)  and  (not A234) );
 a53717a <=( A266  and  A265 );
 a53718a <=( a53717a  and  a53714a );
 a53721a <=( (not A268)  and  (not A267) );
 a53725a <=( (not A301)  and  (not A299) );
 a53726a <=( (not A298)  and  a53725a );
 a53727a <=( a53726a  and  a53721a );
 a53728a <=( a53727a  and  a53718a );
 a53731a <=( (not A167)  and  A170 );
 a53734a <=( (not A199)  and  A166 );
 a53735a <=( a53734a  and  a53731a );
 a53738a <=( (not A202)  and  (not A200) );
 a53741a <=( A233  and  A232 );
 a53742a <=( a53741a  and  a53738a );
 a53743a <=( a53742a  and  a53735a );
 a53746a <=( (not A235)  and  (not A234) );
 a53749a <=( (not A266)  and  (not A265) );
 a53750a <=( a53749a  and  a53746a );
 a53753a <=( A298  and  (not A268) );
 a53757a <=( (not A301)  and  (not A300) );
 a53758a <=( A299  and  a53757a );
 a53759a <=( a53758a  and  a53753a );
 a53760a <=( a53759a  and  a53750a );
 a53763a <=( (not A167)  and  A170 );
 a53766a <=( (not A199)  and  A166 );
 a53767a <=( a53766a  and  a53763a );
 a53770a <=( (not A202)  and  (not A200) );
 a53773a <=( (not A233)  and  (not A232) );
 a53774a <=( a53773a  and  a53770a );
 a53775a <=( a53774a  and  a53767a );
 a53778a <=( A265  and  (not A235) );
 a53781a <=( (not A267)  and  A266 );
 a53782a <=( a53781a  and  a53778a );
 a53785a <=( A298  and  (not A268) );
 a53789a <=( (not A301)  and  (not A300) );
 a53790a <=( A299  and  a53789a );
 a53791a <=( a53790a  and  a53785a );
 a53792a <=( a53791a  and  a53782a );
 a53795a <=( A199  and  A169 );
 a53798a <=( (not A201)  and  A200 );
 a53799a <=( a53798a  and  a53795a );
 a53802a <=( A232  and  (not A202) );
 a53805a <=( (not A234)  and  A233 );
 a53806a <=( a53805a  and  a53802a );
 a53807a <=( a53806a  and  a53799a );
 a53810a <=( A265  and  (not A235) );
 a53813a <=( (not A267)  and  A266 );
 a53814a <=( a53813a  and  a53810a );
 a53817a <=( A298  and  (not A268) );
 a53821a <=( (not A301)  and  (not A300) );
 a53822a <=( A299  and  a53821a );
 a53823a <=( a53822a  and  a53817a );
 a53824a <=( a53823a  and  a53814a );
 a53827a <=( (not A167)  and  (not A169) );
 a53830a <=( A199  and  (not A166) );
 a53831a <=( a53830a  and  a53827a );
 a53834a <=( A232  and  A201 );
 a53837a <=( (not A234)  and  A233 );
 a53838a <=( a53837a  and  a53834a );
 a53839a <=( a53838a  and  a53831a );
 a53842a <=( A265  and  (not A235) );
 a53845a <=( (not A267)  and  A266 );
 a53846a <=( a53845a  and  a53842a );
 a53849a <=( A298  and  (not A268) );
 a53853a <=( (not A301)  and  (not A300) );
 a53854a <=( A299  and  a53853a );
 a53855a <=( a53854a  and  a53849a );
 a53856a <=( a53855a  and  a53846a );
 a53859a <=( (not A167)  and  (not A169) );
 a53862a <=( A200  and  (not A166) );
 a53863a <=( a53862a  and  a53859a );
 a53866a <=( A232  and  A201 );
 a53869a <=( (not A234)  and  A233 );
 a53870a <=( a53869a  and  a53866a );
 a53871a <=( a53870a  and  a53863a );
 a53874a <=( A265  and  (not A235) );
 a53877a <=( (not A267)  and  A266 );
 a53878a <=( a53877a  and  a53874a );
 a53881a <=( A298  and  (not A268) );
 a53885a <=( (not A301)  and  (not A300) );
 a53886a <=( A299  and  a53885a );
 a53887a <=( a53886a  and  a53881a );
 a53888a <=( a53887a  and  a53878a );
 a53891a <=( (not A167)  and  (not A169) );
 a53894a <=( (not A199)  and  (not A166) );
 a53895a <=( a53894a  and  a53891a );
 a53898a <=( A203  and  A200 );
 a53901a <=( (not A235)  and  (not A234) );
 a53902a <=( a53901a  and  a53898a );
 a53903a <=( a53902a  and  a53895a );
 a53906a <=( A265  and  (not A236) );
 a53909a <=( (not A267)  and  A266 );
 a53910a <=( a53909a  and  a53906a );
 a53913a <=( A298  and  (not A268) );
 a53917a <=( (not A301)  and  (not A300) );
 a53918a <=( A299  and  a53917a );
 a53919a <=( a53918a  and  a53913a );
 a53920a <=( a53919a  and  a53910a );
 a53923a <=( (not A167)  and  (not A169) );
 a53926a <=( (not A199)  and  (not A166) );
 a53927a <=( a53926a  and  a53923a );
 a53930a <=( A203  and  A200 );
 a53933a <=( A233  and  A232 );
 a53934a <=( a53933a  and  a53930a );
 a53935a <=( a53934a  and  a53927a );
 a53938a <=( (not A235)  and  (not A234) );
 a53941a <=( (not A268)  and  (not A267) );
 a53942a <=( a53941a  and  a53938a );
 a53945a <=( A298  and  (not A269) );
 a53949a <=( (not A301)  and  (not A300) );
 a53950a <=( A299  and  a53949a );
 a53951a <=( a53950a  and  a53945a );
 a53952a <=( a53951a  and  a53942a );
 a53955a <=( (not A167)  and  (not A169) );
 a53958a <=( (not A199)  and  (not A166) );
 a53959a <=( a53958a  and  a53955a );
 a53962a <=( A203  and  A200 );
 a53965a <=( A233  and  A232 );
 a53966a <=( a53965a  and  a53962a );
 a53967a <=( a53966a  and  a53959a );
 a53970a <=( (not A235)  and  (not A234) );
 a53973a <=( A266  and  A265 );
 a53974a <=( a53973a  and  a53970a );
 a53977a <=( (not A268)  and  (not A267) );
 a53981a <=( (not A302)  and  (not A301) );
 a53982a <=( (not A300)  and  a53981a );
 a53983a <=( a53982a  and  a53977a );
 a53984a <=( a53983a  and  a53974a );
 a53987a <=( (not A167)  and  (not A169) );
 a53990a <=( (not A199)  and  (not A166) );
 a53991a <=( a53990a  and  a53987a );
 a53994a <=( A203  and  A200 );
 a53997a <=( A233  and  A232 );
 a53998a <=( a53997a  and  a53994a );
 a53999a <=( a53998a  and  a53991a );
 a54002a <=( (not A235)  and  (not A234) );
 a54005a <=( A266  and  A265 );
 a54006a <=( a54005a  and  a54002a );
 a54009a <=( (not A268)  and  (not A267) );
 a54013a <=( (not A301)  and  (not A299) );
 a54014a <=( (not A298)  and  a54013a );
 a54015a <=( a54014a  and  a54009a );
 a54016a <=( a54015a  and  a54006a );
 a54019a <=( (not A167)  and  (not A169) );
 a54022a <=( (not A199)  and  (not A166) );
 a54023a <=( a54022a  and  a54019a );
 a54026a <=( A203  and  A200 );
 a54029a <=( A233  and  A232 );
 a54030a <=( a54029a  and  a54026a );
 a54031a <=( a54030a  and  a54023a );
 a54034a <=( (not A235)  and  (not A234) );
 a54037a <=( (not A266)  and  (not A265) );
 a54038a <=( a54037a  and  a54034a );
 a54041a <=( A298  and  (not A268) );
 a54045a <=( (not A301)  and  (not A300) );
 a54046a <=( A299  and  a54045a );
 a54047a <=( a54046a  and  a54041a );
 a54048a <=( a54047a  and  a54038a );
 a54051a <=( (not A167)  and  (not A169) );
 a54054a <=( (not A199)  and  (not A166) );
 a54055a <=( a54054a  and  a54051a );
 a54058a <=( A203  and  A200 );
 a54061a <=( (not A233)  and  (not A232) );
 a54062a <=( a54061a  and  a54058a );
 a54063a <=( a54062a  and  a54055a );
 a54066a <=( A265  and  (not A235) );
 a54069a <=( (not A267)  and  A266 );
 a54070a <=( a54069a  and  a54066a );
 a54073a <=( A298  and  (not A268) );
 a54077a <=( (not A301)  and  (not A300) );
 a54078a <=( A299  and  a54077a );
 a54079a <=( a54078a  and  a54073a );
 a54080a <=( a54079a  and  a54070a );
 a54083a <=( (not A167)  and  (not A169) );
 a54086a <=( A199  and  (not A166) );
 a54087a <=( a54086a  and  a54083a );
 a54090a <=( A203  and  (not A200) );
 a54093a <=( (not A235)  and  (not A234) );
 a54094a <=( a54093a  and  a54090a );
 a54095a <=( a54094a  and  a54087a );
 a54098a <=( A265  and  (not A236) );
 a54101a <=( (not A267)  and  A266 );
 a54102a <=( a54101a  and  a54098a );
 a54105a <=( A298  and  (not A268) );
 a54109a <=( (not A301)  and  (not A300) );
 a54110a <=( A299  and  a54109a );
 a54111a <=( a54110a  and  a54105a );
 a54112a <=( a54111a  and  a54102a );
 a54115a <=( (not A167)  and  (not A169) );
 a54118a <=( A199  and  (not A166) );
 a54119a <=( a54118a  and  a54115a );
 a54122a <=( A203  and  (not A200) );
 a54125a <=( A233  and  A232 );
 a54126a <=( a54125a  and  a54122a );
 a54127a <=( a54126a  and  a54119a );
 a54130a <=( (not A235)  and  (not A234) );
 a54133a <=( (not A268)  and  (not A267) );
 a54134a <=( a54133a  and  a54130a );
 a54137a <=( A298  and  (not A269) );
 a54141a <=( (not A301)  and  (not A300) );
 a54142a <=( A299  and  a54141a );
 a54143a <=( a54142a  and  a54137a );
 a54144a <=( a54143a  and  a54134a );
 a54147a <=( (not A167)  and  (not A169) );
 a54150a <=( A199  and  (not A166) );
 a54151a <=( a54150a  and  a54147a );
 a54154a <=( A203  and  (not A200) );
 a54157a <=( A233  and  A232 );
 a54158a <=( a54157a  and  a54154a );
 a54159a <=( a54158a  and  a54151a );
 a54162a <=( (not A235)  and  (not A234) );
 a54165a <=( A266  and  A265 );
 a54166a <=( a54165a  and  a54162a );
 a54169a <=( (not A268)  and  (not A267) );
 a54173a <=( (not A302)  and  (not A301) );
 a54174a <=( (not A300)  and  a54173a );
 a54175a <=( a54174a  and  a54169a );
 a54176a <=( a54175a  and  a54166a );
 a54179a <=( (not A167)  and  (not A169) );
 a54182a <=( A199  and  (not A166) );
 a54183a <=( a54182a  and  a54179a );
 a54186a <=( A203  and  (not A200) );
 a54189a <=( A233  and  A232 );
 a54190a <=( a54189a  and  a54186a );
 a54191a <=( a54190a  and  a54183a );
 a54194a <=( (not A235)  and  (not A234) );
 a54197a <=( A266  and  A265 );
 a54198a <=( a54197a  and  a54194a );
 a54201a <=( (not A268)  and  (not A267) );
 a54205a <=( (not A301)  and  (not A299) );
 a54206a <=( (not A298)  and  a54205a );
 a54207a <=( a54206a  and  a54201a );
 a54208a <=( a54207a  and  a54198a );
 a54211a <=( (not A167)  and  (not A169) );
 a54214a <=( A199  and  (not A166) );
 a54215a <=( a54214a  and  a54211a );
 a54218a <=( A203  and  (not A200) );
 a54221a <=( A233  and  A232 );
 a54222a <=( a54221a  and  a54218a );
 a54223a <=( a54222a  and  a54215a );
 a54226a <=( (not A235)  and  (not A234) );
 a54229a <=( (not A266)  and  (not A265) );
 a54230a <=( a54229a  and  a54226a );
 a54233a <=( A298  and  (not A268) );
 a54237a <=( (not A301)  and  (not A300) );
 a54238a <=( A299  and  a54237a );
 a54239a <=( a54238a  and  a54233a );
 a54240a <=( a54239a  and  a54230a );
 a54243a <=( (not A167)  and  (not A169) );
 a54246a <=( A199  and  (not A166) );
 a54247a <=( a54246a  and  a54243a );
 a54250a <=( A203  and  (not A200) );
 a54253a <=( (not A233)  and  (not A232) );
 a54254a <=( a54253a  and  a54250a );
 a54255a <=( a54254a  and  a54247a );
 a54258a <=( A265  and  (not A235) );
 a54261a <=( (not A267)  and  A266 );
 a54262a <=( a54261a  and  a54258a );
 a54265a <=( A298  and  (not A268) );
 a54269a <=( (not A301)  and  (not A300) );
 a54270a <=( A299  and  a54269a );
 a54271a <=( a54270a  and  a54265a );
 a54272a <=( a54271a  and  a54262a );
 a54275a <=( (not A168)  and  (not A169) );
 a54278a <=( A166  and  A167 );
 a54279a <=( a54278a  and  a54275a );
 a54282a <=( A232  and  A202 );
 a54285a <=( (not A234)  and  A233 );
 a54286a <=( a54285a  and  a54282a );
 a54287a <=( a54286a  and  a54279a );
 a54290a <=( A265  and  (not A235) );
 a54293a <=( (not A267)  and  A266 );
 a54294a <=( a54293a  and  a54290a );
 a54297a <=( A298  and  (not A268) );
 a54301a <=( (not A301)  and  (not A300) );
 a54302a <=( A299  and  a54301a );
 a54303a <=( a54302a  and  a54297a );
 a54304a <=( a54303a  and  a54294a );
 a54307a <=( (not A168)  and  (not A169) );
 a54310a <=( A166  and  A167 );
 a54311a <=( a54310a  and  a54307a );
 a54314a <=( A201  and  A199 );
 a54317a <=( (not A235)  and  (not A234) );
 a54318a <=( a54317a  and  a54314a );
 a54319a <=( a54318a  and  a54311a );
 a54322a <=( A265  and  (not A236) );
 a54325a <=( (not A267)  and  A266 );
 a54326a <=( a54325a  and  a54322a );
 a54329a <=( A298  and  (not A268) );
 a54333a <=( (not A301)  and  (not A300) );
 a54334a <=( A299  and  a54333a );
 a54335a <=( a54334a  and  a54329a );
 a54336a <=( a54335a  and  a54326a );
 a54339a <=( (not A168)  and  (not A169) );
 a54342a <=( A166  and  A167 );
 a54343a <=( a54342a  and  a54339a );
 a54346a <=( A201  and  A199 );
 a54349a <=( A233  and  A232 );
 a54350a <=( a54349a  and  a54346a );
 a54351a <=( a54350a  and  a54343a );
 a54354a <=( (not A235)  and  (not A234) );
 a54357a <=( (not A268)  and  (not A267) );
 a54358a <=( a54357a  and  a54354a );
 a54361a <=( A298  and  (not A269) );
 a54365a <=( (not A301)  and  (not A300) );
 a54366a <=( A299  and  a54365a );
 a54367a <=( a54366a  and  a54361a );
 a54368a <=( a54367a  and  a54358a );
 a54371a <=( (not A168)  and  (not A169) );
 a54374a <=( A166  and  A167 );
 a54375a <=( a54374a  and  a54371a );
 a54378a <=( A201  and  A199 );
 a54381a <=( A233  and  A232 );
 a54382a <=( a54381a  and  a54378a );
 a54383a <=( a54382a  and  a54375a );
 a54386a <=( (not A235)  and  (not A234) );
 a54389a <=( A266  and  A265 );
 a54390a <=( a54389a  and  a54386a );
 a54393a <=( (not A268)  and  (not A267) );
 a54397a <=( (not A302)  and  (not A301) );
 a54398a <=( (not A300)  and  a54397a );
 a54399a <=( a54398a  and  a54393a );
 a54400a <=( a54399a  and  a54390a );
 a54403a <=( (not A168)  and  (not A169) );
 a54406a <=( A166  and  A167 );
 a54407a <=( a54406a  and  a54403a );
 a54410a <=( A201  and  A199 );
 a54413a <=( A233  and  A232 );
 a54414a <=( a54413a  and  a54410a );
 a54415a <=( a54414a  and  a54407a );
 a54418a <=( (not A235)  and  (not A234) );
 a54421a <=( A266  and  A265 );
 a54422a <=( a54421a  and  a54418a );
 a54425a <=( (not A268)  and  (not A267) );
 a54429a <=( (not A301)  and  (not A299) );
 a54430a <=( (not A298)  and  a54429a );
 a54431a <=( a54430a  and  a54425a );
 a54432a <=( a54431a  and  a54422a );
 a54435a <=( (not A168)  and  (not A169) );
 a54438a <=( A166  and  A167 );
 a54439a <=( a54438a  and  a54435a );
 a54442a <=( A201  and  A199 );
 a54445a <=( A233  and  A232 );
 a54446a <=( a54445a  and  a54442a );
 a54447a <=( a54446a  and  a54439a );
 a54450a <=( (not A235)  and  (not A234) );
 a54453a <=( (not A266)  and  (not A265) );
 a54454a <=( a54453a  and  a54450a );
 a54457a <=( A298  and  (not A268) );
 a54461a <=( (not A301)  and  (not A300) );
 a54462a <=( A299  and  a54461a );
 a54463a <=( a54462a  and  a54457a );
 a54464a <=( a54463a  and  a54454a );
 a54467a <=( (not A168)  and  (not A169) );
 a54470a <=( A166  and  A167 );
 a54471a <=( a54470a  and  a54467a );
 a54474a <=( A201  and  A199 );
 a54477a <=( (not A233)  and  (not A232) );
 a54478a <=( a54477a  and  a54474a );
 a54479a <=( a54478a  and  a54471a );
 a54482a <=( A265  and  (not A235) );
 a54485a <=( (not A267)  and  A266 );
 a54486a <=( a54485a  and  a54482a );
 a54489a <=( A298  and  (not A268) );
 a54493a <=( (not A301)  and  (not A300) );
 a54494a <=( A299  and  a54493a );
 a54495a <=( a54494a  and  a54489a );
 a54496a <=( a54495a  and  a54486a );
 a54499a <=( (not A168)  and  (not A169) );
 a54502a <=( A166  and  A167 );
 a54503a <=( a54502a  and  a54499a );
 a54506a <=( A201  and  A200 );
 a54509a <=( (not A235)  and  (not A234) );
 a54510a <=( a54509a  and  a54506a );
 a54511a <=( a54510a  and  a54503a );
 a54514a <=( A265  and  (not A236) );
 a54517a <=( (not A267)  and  A266 );
 a54518a <=( a54517a  and  a54514a );
 a54521a <=( A298  and  (not A268) );
 a54525a <=( (not A301)  and  (not A300) );
 a54526a <=( A299  and  a54525a );
 a54527a <=( a54526a  and  a54521a );
 a54528a <=( a54527a  and  a54518a );
 a54531a <=( (not A168)  and  (not A169) );
 a54534a <=( A166  and  A167 );
 a54535a <=( a54534a  and  a54531a );
 a54538a <=( A201  and  A200 );
 a54541a <=( A233  and  A232 );
 a54542a <=( a54541a  and  a54538a );
 a54543a <=( a54542a  and  a54535a );
 a54546a <=( (not A235)  and  (not A234) );
 a54549a <=( (not A268)  and  (not A267) );
 a54550a <=( a54549a  and  a54546a );
 a54553a <=( A298  and  (not A269) );
 a54557a <=( (not A301)  and  (not A300) );
 a54558a <=( A299  and  a54557a );
 a54559a <=( a54558a  and  a54553a );
 a54560a <=( a54559a  and  a54550a );
 a54563a <=( (not A168)  and  (not A169) );
 a54566a <=( A166  and  A167 );
 a54567a <=( a54566a  and  a54563a );
 a54570a <=( A201  and  A200 );
 a54573a <=( A233  and  A232 );
 a54574a <=( a54573a  and  a54570a );
 a54575a <=( a54574a  and  a54567a );
 a54578a <=( (not A235)  and  (not A234) );
 a54581a <=( A266  and  A265 );
 a54582a <=( a54581a  and  a54578a );
 a54585a <=( (not A268)  and  (not A267) );
 a54589a <=( (not A302)  and  (not A301) );
 a54590a <=( (not A300)  and  a54589a );
 a54591a <=( a54590a  and  a54585a );
 a54592a <=( a54591a  and  a54582a );
 a54595a <=( (not A168)  and  (not A169) );
 a54598a <=( A166  and  A167 );
 a54599a <=( a54598a  and  a54595a );
 a54602a <=( A201  and  A200 );
 a54605a <=( A233  and  A232 );
 a54606a <=( a54605a  and  a54602a );
 a54607a <=( a54606a  and  a54599a );
 a54610a <=( (not A235)  and  (not A234) );
 a54613a <=( A266  and  A265 );
 a54614a <=( a54613a  and  a54610a );
 a54617a <=( (not A268)  and  (not A267) );
 a54621a <=( (not A301)  and  (not A299) );
 a54622a <=( (not A298)  and  a54621a );
 a54623a <=( a54622a  and  a54617a );
 a54624a <=( a54623a  and  a54614a );
 a54627a <=( (not A168)  and  (not A169) );
 a54630a <=( A166  and  A167 );
 a54631a <=( a54630a  and  a54627a );
 a54634a <=( A201  and  A200 );
 a54637a <=( A233  and  A232 );
 a54638a <=( a54637a  and  a54634a );
 a54639a <=( a54638a  and  a54631a );
 a54642a <=( (not A235)  and  (not A234) );
 a54645a <=( (not A266)  and  (not A265) );
 a54646a <=( a54645a  and  a54642a );
 a54649a <=( A298  and  (not A268) );
 a54653a <=( (not A301)  and  (not A300) );
 a54654a <=( A299  and  a54653a );
 a54655a <=( a54654a  and  a54649a );
 a54656a <=( a54655a  and  a54646a );
 a54659a <=( (not A168)  and  (not A169) );
 a54662a <=( A166  and  A167 );
 a54663a <=( a54662a  and  a54659a );
 a54666a <=( A201  and  A200 );
 a54669a <=( (not A233)  and  (not A232) );
 a54670a <=( a54669a  and  a54666a );
 a54671a <=( a54670a  and  a54663a );
 a54674a <=( A265  and  (not A235) );
 a54677a <=( (not A267)  and  A266 );
 a54678a <=( a54677a  and  a54674a );
 a54681a <=( A298  and  (not A268) );
 a54685a <=( (not A301)  and  (not A300) );
 a54686a <=( A299  and  a54685a );
 a54687a <=( a54686a  and  a54681a );
 a54688a <=( a54687a  and  a54678a );
 a54691a <=( (not A168)  and  (not A169) );
 a54694a <=( A166  and  A167 );
 a54695a <=( a54694a  and  a54691a );
 a54698a <=( A200  and  (not A199) );
 a54701a <=( (not A234)  and  A203 );
 a54702a <=( a54701a  and  a54698a );
 a54703a <=( a54702a  and  a54695a );
 a54706a <=( (not A236)  and  (not A235) );
 a54709a <=( (not A268)  and  (not A267) );
 a54710a <=( a54709a  and  a54706a );
 a54713a <=( A298  and  (not A269) );
 a54717a <=( (not A301)  and  (not A300) );
 a54718a <=( A299  and  a54717a );
 a54719a <=( a54718a  and  a54713a );
 a54720a <=( a54719a  and  a54710a );
 a54723a <=( (not A168)  and  (not A169) );
 a54726a <=( A166  and  A167 );
 a54727a <=( a54726a  and  a54723a );
 a54730a <=( A200  and  (not A199) );
 a54733a <=( (not A234)  and  A203 );
 a54734a <=( a54733a  and  a54730a );
 a54735a <=( a54734a  and  a54727a );
 a54738a <=( (not A236)  and  (not A235) );
 a54741a <=( A266  and  A265 );
 a54742a <=( a54741a  and  a54738a );
 a54745a <=( (not A268)  and  (not A267) );
 a54749a <=( (not A302)  and  (not A301) );
 a54750a <=( (not A300)  and  a54749a );
 a54751a <=( a54750a  and  a54745a );
 a54752a <=( a54751a  and  a54742a );
 a54755a <=( (not A168)  and  (not A169) );
 a54758a <=( A166  and  A167 );
 a54759a <=( a54758a  and  a54755a );
 a54762a <=( A200  and  (not A199) );
 a54765a <=( (not A234)  and  A203 );
 a54766a <=( a54765a  and  a54762a );
 a54767a <=( a54766a  and  a54759a );
 a54770a <=( (not A236)  and  (not A235) );
 a54773a <=( A266  and  A265 );
 a54774a <=( a54773a  and  a54770a );
 a54777a <=( (not A268)  and  (not A267) );
 a54781a <=( (not A301)  and  (not A299) );
 a54782a <=( (not A298)  and  a54781a );
 a54783a <=( a54782a  and  a54777a );
 a54784a <=( a54783a  and  a54774a );
 a54787a <=( (not A168)  and  (not A169) );
 a54790a <=( A166  and  A167 );
 a54791a <=( a54790a  and  a54787a );
 a54794a <=( A200  and  (not A199) );
 a54797a <=( (not A234)  and  A203 );
 a54798a <=( a54797a  and  a54794a );
 a54799a <=( a54798a  and  a54791a );
 a54802a <=( (not A236)  and  (not A235) );
 a54805a <=( (not A266)  and  (not A265) );
 a54806a <=( a54805a  and  a54802a );
 a54809a <=( A298  and  (not A268) );
 a54813a <=( (not A301)  and  (not A300) );
 a54814a <=( A299  and  a54813a );
 a54815a <=( a54814a  and  a54809a );
 a54816a <=( a54815a  and  a54806a );
 a54819a <=( (not A168)  and  (not A169) );
 a54822a <=( A166  and  A167 );
 a54823a <=( a54822a  and  a54819a );
 a54826a <=( A200  and  (not A199) );
 a54829a <=( A232  and  A203 );
 a54830a <=( a54829a  and  a54826a );
 a54831a <=( a54830a  and  a54823a );
 a54834a <=( (not A234)  and  A233 );
 a54837a <=( (not A267)  and  (not A235) );
 a54838a <=( a54837a  and  a54834a );
 a54841a <=( (not A269)  and  (not A268) );
 a54845a <=( (not A302)  and  (not A301) );
 a54846a <=( (not A300)  and  a54845a );
 a54847a <=( a54846a  and  a54841a );
 a54848a <=( a54847a  and  a54838a );
 a54851a <=( (not A168)  and  (not A169) );
 a54854a <=( A166  and  A167 );
 a54855a <=( a54854a  and  a54851a );
 a54858a <=( A200  and  (not A199) );
 a54861a <=( A232  and  A203 );
 a54862a <=( a54861a  and  a54858a );
 a54863a <=( a54862a  and  a54855a );
 a54866a <=( (not A234)  and  A233 );
 a54869a <=( (not A267)  and  (not A235) );
 a54870a <=( a54869a  and  a54866a );
 a54873a <=( (not A269)  and  (not A268) );
 a54877a <=( (not A301)  and  (not A299) );
 a54878a <=( (not A298)  and  a54877a );
 a54879a <=( a54878a  and  a54873a );
 a54880a <=( a54879a  and  a54870a );
 a54883a <=( (not A168)  and  (not A169) );
 a54886a <=( A166  and  A167 );
 a54887a <=( a54886a  and  a54883a );
 a54890a <=( A200  and  (not A199) );
 a54893a <=( A232  and  A203 );
 a54894a <=( a54893a  and  a54890a );
 a54895a <=( a54894a  and  a54887a );
 a54898a <=( (not A234)  and  A233 );
 a54901a <=( (not A265)  and  (not A235) );
 a54902a <=( a54901a  and  a54898a );
 a54905a <=( (not A268)  and  (not A266) );
 a54909a <=( (not A302)  and  (not A301) );
 a54910a <=( (not A300)  and  a54909a );
 a54911a <=( a54910a  and  a54905a );
 a54912a <=( a54911a  and  a54902a );
 a54915a <=( (not A168)  and  (not A169) );
 a54918a <=( A166  and  A167 );
 a54919a <=( a54918a  and  a54915a );
 a54922a <=( A200  and  (not A199) );
 a54925a <=( A232  and  A203 );
 a54926a <=( a54925a  and  a54922a );
 a54927a <=( a54926a  and  a54919a );
 a54930a <=( (not A234)  and  A233 );
 a54933a <=( (not A265)  and  (not A235) );
 a54934a <=( a54933a  and  a54930a );
 a54937a <=( (not A268)  and  (not A266) );
 a54941a <=( (not A301)  and  (not A299) );
 a54942a <=( (not A298)  and  a54941a );
 a54943a <=( a54942a  and  a54937a );
 a54944a <=( a54943a  and  a54934a );
 a54947a <=( (not A168)  and  (not A169) );
 a54950a <=( A166  and  A167 );
 a54951a <=( a54950a  and  a54947a );
 a54954a <=( A200  and  (not A199) );
 a54957a <=( (not A232)  and  A203 );
 a54958a <=( a54957a  and  a54954a );
 a54959a <=( a54958a  and  a54951a );
 a54962a <=( (not A235)  and  (not A233) );
 a54965a <=( (not A268)  and  (not A267) );
 a54966a <=( a54965a  and  a54962a );
 a54969a <=( A298  and  (not A269) );
 a54973a <=( (not A301)  and  (not A300) );
 a54974a <=( A299  and  a54973a );
 a54975a <=( a54974a  and  a54969a );
 a54976a <=( a54975a  and  a54966a );
 a54979a <=( (not A168)  and  (not A169) );
 a54982a <=( A166  and  A167 );
 a54983a <=( a54982a  and  a54979a );
 a54986a <=( A200  and  (not A199) );
 a54989a <=( (not A232)  and  A203 );
 a54990a <=( a54989a  and  a54986a );
 a54991a <=( a54990a  and  a54983a );
 a54994a <=( (not A235)  and  (not A233) );
 a54997a <=( A266  and  A265 );
 a54998a <=( a54997a  and  a54994a );
 a55001a <=( (not A268)  and  (not A267) );
 a55005a <=( (not A302)  and  (not A301) );
 a55006a <=( (not A300)  and  a55005a );
 a55007a <=( a55006a  and  a55001a );
 a55008a <=( a55007a  and  a54998a );
 a55011a <=( (not A168)  and  (not A169) );
 a55014a <=( A166  and  A167 );
 a55015a <=( a55014a  and  a55011a );
 a55018a <=( A200  and  (not A199) );
 a55021a <=( (not A232)  and  A203 );
 a55022a <=( a55021a  and  a55018a );
 a55023a <=( a55022a  and  a55015a );
 a55026a <=( (not A235)  and  (not A233) );
 a55029a <=( A266  and  A265 );
 a55030a <=( a55029a  and  a55026a );
 a55033a <=( (not A268)  and  (not A267) );
 a55037a <=( (not A301)  and  (not A299) );
 a55038a <=( (not A298)  and  a55037a );
 a55039a <=( a55038a  and  a55033a );
 a55040a <=( a55039a  and  a55030a );
 a55043a <=( (not A168)  and  (not A169) );
 a55046a <=( A166  and  A167 );
 a55047a <=( a55046a  and  a55043a );
 a55050a <=( A200  and  (not A199) );
 a55053a <=( (not A232)  and  A203 );
 a55054a <=( a55053a  and  a55050a );
 a55055a <=( a55054a  and  a55047a );
 a55058a <=( (not A235)  and  (not A233) );
 a55061a <=( (not A266)  and  (not A265) );
 a55062a <=( a55061a  and  a55058a );
 a55065a <=( A298  and  (not A268) );
 a55069a <=( (not A301)  and  (not A300) );
 a55070a <=( A299  and  a55069a );
 a55071a <=( a55070a  and  a55065a );
 a55072a <=( a55071a  and  a55062a );
 a55075a <=( (not A168)  and  (not A169) );
 a55078a <=( A166  and  A167 );
 a55079a <=( a55078a  and  a55075a );
 a55082a <=( (not A200)  and  A199 );
 a55085a <=( (not A234)  and  A203 );
 a55086a <=( a55085a  and  a55082a );
 a55087a <=( a55086a  and  a55079a );
 a55090a <=( (not A236)  and  (not A235) );
 a55093a <=( (not A268)  and  (not A267) );
 a55094a <=( a55093a  and  a55090a );
 a55097a <=( A298  and  (not A269) );
 a55101a <=( (not A301)  and  (not A300) );
 a55102a <=( A299  and  a55101a );
 a55103a <=( a55102a  and  a55097a );
 a55104a <=( a55103a  and  a55094a );
 a55107a <=( (not A168)  and  (not A169) );
 a55110a <=( A166  and  A167 );
 a55111a <=( a55110a  and  a55107a );
 a55114a <=( (not A200)  and  A199 );
 a55117a <=( (not A234)  and  A203 );
 a55118a <=( a55117a  and  a55114a );
 a55119a <=( a55118a  and  a55111a );
 a55122a <=( (not A236)  and  (not A235) );
 a55125a <=( A266  and  A265 );
 a55126a <=( a55125a  and  a55122a );
 a55129a <=( (not A268)  and  (not A267) );
 a55133a <=( (not A302)  and  (not A301) );
 a55134a <=( (not A300)  and  a55133a );
 a55135a <=( a55134a  and  a55129a );
 a55136a <=( a55135a  and  a55126a );
 a55139a <=( (not A168)  and  (not A169) );
 a55142a <=( A166  and  A167 );
 a55143a <=( a55142a  and  a55139a );
 a55146a <=( (not A200)  and  A199 );
 a55149a <=( (not A234)  and  A203 );
 a55150a <=( a55149a  and  a55146a );
 a55151a <=( a55150a  and  a55143a );
 a55154a <=( (not A236)  and  (not A235) );
 a55157a <=( A266  and  A265 );
 a55158a <=( a55157a  and  a55154a );
 a55161a <=( (not A268)  and  (not A267) );
 a55165a <=( (not A301)  and  (not A299) );
 a55166a <=( (not A298)  and  a55165a );
 a55167a <=( a55166a  and  a55161a );
 a55168a <=( a55167a  and  a55158a );
 a55171a <=( (not A168)  and  (not A169) );
 a55174a <=( A166  and  A167 );
 a55175a <=( a55174a  and  a55171a );
 a55178a <=( (not A200)  and  A199 );
 a55181a <=( (not A234)  and  A203 );
 a55182a <=( a55181a  and  a55178a );
 a55183a <=( a55182a  and  a55175a );
 a55186a <=( (not A236)  and  (not A235) );
 a55189a <=( (not A266)  and  (not A265) );
 a55190a <=( a55189a  and  a55186a );
 a55193a <=( A298  and  (not A268) );
 a55197a <=( (not A301)  and  (not A300) );
 a55198a <=( A299  and  a55197a );
 a55199a <=( a55198a  and  a55193a );
 a55200a <=( a55199a  and  a55190a );
 a55203a <=( (not A168)  and  (not A169) );
 a55206a <=( A166  and  A167 );
 a55207a <=( a55206a  and  a55203a );
 a55210a <=( (not A200)  and  A199 );
 a55213a <=( A232  and  A203 );
 a55214a <=( a55213a  and  a55210a );
 a55215a <=( a55214a  and  a55207a );
 a55218a <=( (not A234)  and  A233 );
 a55221a <=( (not A267)  and  (not A235) );
 a55222a <=( a55221a  and  a55218a );
 a55225a <=( (not A269)  and  (not A268) );
 a55229a <=( (not A302)  and  (not A301) );
 a55230a <=( (not A300)  and  a55229a );
 a55231a <=( a55230a  and  a55225a );
 a55232a <=( a55231a  and  a55222a );
 a55235a <=( (not A168)  and  (not A169) );
 a55238a <=( A166  and  A167 );
 a55239a <=( a55238a  and  a55235a );
 a55242a <=( (not A200)  and  A199 );
 a55245a <=( A232  and  A203 );
 a55246a <=( a55245a  and  a55242a );
 a55247a <=( a55246a  and  a55239a );
 a55250a <=( (not A234)  and  A233 );
 a55253a <=( (not A267)  and  (not A235) );
 a55254a <=( a55253a  and  a55250a );
 a55257a <=( (not A269)  and  (not A268) );
 a55261a <=( (not A301)  and  (not A299) );
 a55262a <=( (not A298)  and  a55261a );
 a55263a <=( a55262a  and  a55257a );
 a55264a <=( a55263a  and  a55254a );
 a55267a <=( (not A168)  and  (not A169) );
 a55270a <=( A166  and  A167 );
 a55271a <=( a55270a  and  a55267a );
 a55274a <=( (not A200)  and  A199 );
 a55277a <=( A232  and  A203 );
 a55278a <=( a55277a  and  a55274a );
 a55279a <=( a55278a  and  a55271a );
 a55282a <=( (not A234)  and  A233 );
 a55285a <=( (not A265)  and  (not A235) );
 a55286a <=( a55285a  and  a55282a );
 a55289a <=( (not A268)  and  (not A266) );
 a55293a <=( (not A302)  and  (not A301) );
 a55294a <=( (not A300)  and  a55293a );
 a55295a <=( a55294a  and  a55289a );
 a55296a <=( a55295a  and  a55286a );
 a55299a <=( (not A168)  and  (not A169) );
 a55302a <=( A166  and  A167 );
 a55303a <=( a55302a  and  a55299a );
 a55306a <=( (not A200)  and  A199 );
 a55309a <=( A232  and  A203 );
 a55310a <=( a55309a  and  a55306a );
 a55311a <=( a55310a  and  a55303a );
 a55314a <=( (not A234)  and  A233 );
 a55317a <=( (not A265)  and  (not A235) );
 a55318a <=( a55317a  and  a55314a );
 a55321a <=( (not A268)  and  (not A266) );
 a55325a <=( (not A301)  and  (not A299) );
 a55326a <=( (not A298)  and  a55325a );
 a55327a <=( a55326a  and  a55321a );
 a55328a <=( a55327a  and  a55318a );
 a55331a <=( (not A168)  and  (not A169) );
 a55334a <=( A166  and  A167 );
 a55335a <=( a55334a  and  a55331a );
 a55338a <=( (not A200)  and  A199 );
 a55341a <=( (not A232)  and  A203 );
 a55342a <=( a55341a  and  a55338a );
 a55343a <=( a55342a  and  a55335a );
 a55346a <=( (not A235)  and  (not A233) );
 a55349a <=( (not A268)  and  (not A267) );
 a55350a <=( a55349a  and  a55346a );
 a55353a <=( A298  and  (not A269) );
 a55357a <=( (not A301)  and  (not A300) );
 a55358a <=( A299  and  a55357a );
 a55359a <=( a55358a  and  a55353a );
 a55360a <=( a55359a  and  a55350a );
 a55363a <=( (not A168)  and  (not A169) );
 a55366a <=( A166  and  A167 );
 a55367a <=( a55366a  and  a55363a );
 a55370a <=( (not A200)  and  A199 );
 a55373a <=( (not A232)  and  A203 );
 a55374a <=( a55373a  and  a55370a );
 a55375a <=( a55374a  and  a55367a );
 a55378a <=( (not A235)  and  (not A233) );
 a55381a <=( A266  and  A265 );
 a55382a <=( a55381a  and  a55378a );
 a55385a <=( (not A268)  and  (not A267) );
 a55389a <=( (not A302)  and  (not A301) );
 a55390a <=( (not A300)  and  a55389a );
 a55391a <=( a55390a  and  a55385a );
 a55392a <=( a55391a  and  a55382a );
 a55395a <=( (not A168)  and  (not A169) );
 a55398a <=( A166  and  A167 );
 a55399a <=( a55398a  and  a55395a );
 a55402a <=( (not A200)  and  A199 );
 a55405a <=( (not A232)  and  A203 );
 a55406a <=( a55405a  and  a55402a );
 a55407a <=( a55406a  and  a55399a );
 a55410a <=( (not A235)  and  (not A233) );
 a55413a <=( A266  and  A265 );
 a55414a <=( a55413a  and  a55410a );
 a55417a <=( (not A268)  and  (not A267) );
 a55421a <=( (not A301)  and  (not A299) );
 a55422a <=( (not A298)  and  a55421a );
 a55423a <=( a55422a  and  a55417a );
 a55424a <=( a55423a  and  a55414a );
 a55427a <=( (not A168)  and  (not A169) );
 a55430a <=( A166  and  A167 );
 a55431a <=( a55430a  and  a55427a );
 a55434a <=( (not A200)  and  A199 );
 a55437a <=( (not A232)  and  A203 );
 a55438a <=( a55437a  and  a55434a );
 a55439a <=( a55438a  and  a55431a );
 a55442a <=( (not A235)  and  (not A233) );
 a55445a <=( (not A266)  and  (not A265) );
 a55446a <=( a55445a  and  a55442a );
 a55449a <=( A298  and  (not A268) );
 a55453a <=( (not A301)  and  (not A300) );
 a55454a <=( A299  and  a55453a );
 a55455a <=( a55454a  and  a55449a );
 a55456a <=( a55455a  and  a55446a );
 a55459a <=( (not A169)  and  (not A170) );
 a55462a <=( A199  and  (not A168) );
 a55463a <=( a55462a  and  a55459a );
 a55466a <=( A232  and  A201 );
 a55469a <=( (not A234)  and  A233 );
 a55470a <=( a55469a  and  a55466a );
 a55471a <=( a55470a  and  a55463a );
 a55474a <=( A265  and  (not A235) );
 a55477a <=( (not A267)  and  A266 );
 a55478a <=( a55477a  and  a55474a );
 a55481a <=( A298  and  (not A268) );
 a55485a <=( (not A301)  and  (not A300) );
 a55486a <=( A299  and  a55485a );
 a55487a <=( a55486a  and  a55481a );
 a55488a <=( a55487a  and  a55478a );
 a55491a <=( (not A169)  and  (not A170) );
 a55494a <=( A200  and  (not A168) );
 a55495a <=( a55494a  and  a55491a );
 a55498a <=( A232  and  A201 );
 a55501a <=( (not A234)  and  A233 );
 a55502a <=( a55501a  and  a55498a );
 a55503a <=( a55502a  and  a55495a );
 a55506a <=( A265  and  (not A235) );
 a55509a <=( (not A267)  and  A266 );
 a55510a <=( a55509a  and  a55506a );
 a55513a <=( A298  and  (not A268) );
 a55517a <=( (not A301)  and  (not A300) );
 a55518a <=( A299  and  a55517a );
 a55519a <=( a55518a  and  a55513a );
 a55520a <=( a55519a  and  a55510a );
 a55523a <=( (not A169)  and  (not A170) );
 a55526a <=( (not A199)  and  (not A168) );
 a55527a <=( a55526a  and  a55523a );
 a55530a <=( A203  and  A200 );
 a55533a <=( (not A235)  and  (not A234) );
 a55534a <=( a55533a  and  a55530a );
 a55535a <=( a55534a  and  a55527a );
 a55538a <=( A265  and  (not A236) );
 a55541a <=( (not A267)  and  A266 );
 a55542a <=( a55541a  and  a55538a );
 a55545a <=( A298  and  (not A268) );
 a55549a <=( (not A301)  and  (not A300) );
 a55550a <=( A299  and  a55549a );
 a55551a <=( a55550a  and  a55545a );
 a55552a <=( a55551a  and  a55542a );
 a55555a <=( (not A169)  and  (not A170) );
 a55558a <=( (not A199)  and  (not A168) );
 a55559a <=( a55558a  and  a55555a );
 a55562a <=( A203  and  A200 );
 a55565a <=( A233  and  A232 );
 a55566a <=( a55565a  and  a55562a );
 a55567a <=( a55566a  and  a55559a );
 a55570a <=( (not A235)  and  (not A234) );
 a55573a <=( (not A268)  and  (not A267) );
 a55574a <=( a55573a  and  a55570a );
 a55577a <=( A298  and  (not A269) );
 a55581a <=( (not A301)  and  (not A300) );
 a55582a <=( A299  and  a55581a );
 a55583a <=( a55582a  and  a55577a );
 a55584a <=( a55583a  and  a55574a );
 a55587a <=( (not A169)  and  (not A170) );
 a55590a <=( (not A199)  and  (not A168) );
 a55591a <=( a55590a  and  a55587a );
 a55594a <=( A203  and  A200 );
 a55597a <=( A233  and  A232 );
 a55598a <=( a55597a  and  a55594a );
 a55599a <=( a55598a  and  a55591a );
 a55602a <=( (not A235)  and  (not A234) );
 a55605a <=( A266  and  A265 );
 a55606a <=( a55605a  and  a55602a );
 a55609a <=( (not A268)  and  (not A267) );
 a55613a <=( (not A302)  and  (not A301) );
 a55614a <=( (not A300)  and  a55613a );
 a55615a <=( a55614a  and  a55609a );
 a55616a <=( a55615a  and  a55606a );
 a55619a <=( (not A169)  and  (not A170) );
 a55622a <=( (not A199)  and  (not A168) );
 a55623a <=( a55622a  and  a55619a );
 a55626a <=( A203  and  A200 );
 a55629a <=( A233  and  A232 );
 a55630a <=( a55629a  and  a55626a );
 a55631a <=( a55630a  and  a55623a );
 a55634a <=( (not A235)  and  (not A234) );
 a55637a <=( A266  and  A265 );
 a55638a <=( a55637a  and  a55634a );
 a55641a <=( (not A268)  and  (not A267) );
 a55645a <=( (not A301)  and  (not A299) );
 a55646a <=( (not A298)  and  a55645a );
 a55647a <=( a55646a  and  a55641a );
 a55648a <=( a55647a  and  a55638a );
 a55651a <=( (not A169)  and  (not A170) );
 a55654a <=( (not A199)  and  (not A168) );
 a55655a <=( a55654a  and  a55651a );
 a55658a <=( A203  and  A200 );
 a55661a <=( A233  and  A232 );
 a55662a <=( a55661a  and  a55658a );
 a55663a <=( a55662a  and  a55655a );
 a55666a <=( (not A235)  and  (not A234) );
 a55669a <=( (not A266)  and  (not A265) );
 a55670a <=( a55669a  and  a55666a );
 a55673a <=( A298  and  (not A268) );
 a55677a <=( (not A301)  and  (not A300) );
 a55678a <=( A299  and  a55677a );
 a55679a <=( a55678a  and  a55673a );
 a55680a <=( a55679a  and  a55670a );
 a55683a <=( (not A169)  and  (not A170) );
 a55686a <=( (not A199)  and  (not A168) );
 a55687a <=( a55686a  and  a55683a );
 a55690a <=( A203  and  A200 );
 a55693a <=( (not A233)  and  (not A232) );
 a55694a <=( a55693a  and  a55690a );
 a55695a <=( a55694a  and  a55687a );
 a55698a <=( A265  and  (not A235) );
 a55701a <=( (not A267)  and  A266 );
 a55702a <=( a55701a  and  a55698a );
 a55705a <=( A298  and  (not A268) );
 a55709a <=( (not A301)  and  (not A300) );
 a55710a <=( A299  and  a55709a );
 a55711a <=( a55710a  and  a55705a );
 a55712a <=( a55711a  and  a55702a );
 a55715a <=( (not A169)  and  (not A170) );
 a55718a <=( A199  and  (not A168) );
 a55719a <=( a55718a  and  a55715a );
 a55722a <=( A203  and  (not A200) );
 a55725a <=( (not A235)  and  (not A234) );
 a55726a <=( a55725a  and  a55722a );
 a55727a <=( a55726a  and  a55719a );
 a55730a <=( A265  and  (not A236) );
 a55733a <=( (not A267)  and  A266 );
 a55734a <=( a55733a  and  a55730a );
 a55737a <=( A298  and  (not A268) );
 a55741a <=( (not A301)  and  (not A300) );
 a55742a <=( A299  and  a55741a );
 a55743a <=( a55742a  and  a55737a );
 a55744a <=( a55743a  and  a55734a );
 a55747a <=( (not A169)  and  (not A170) );
 a55750a <=( A199  and  (not A168) );
 a55751a <=( a55750a  and  a55747a );
 a55754a <=( A203  and  (not A200) );
 a55757a <=( A233  and  A232 );
 a55758a <=( a55757a  and  a55754a );
 a55759a <=( a55758a  and  a55751a );
 a55762a <=( (not A235)  and  (not A234) );
 a55765a <=( (not A268)  and  (not A267) );
 a55766a <=( a55765a  and  a55762a );
 a55769a <=( A298  and  (not A269) );
 a55773a <=( (not A301)  and  (not A300) );
 a55774a <=( A299  and  a55773a );
 a55775a <=( a55774a  and  a55769a );
 a55776a <=( a55775a  and  a55766a );
 a55779a <=( (not A169)  and  (not A170) );
 a55782a <=( A199  and  (not A168) );
 a55783a <=( a55782a  and  a55779a );
 a55786a <=( A203  and  (not A200) );
 a55789a <=( A233  and  A232 );
 a55790a <=( a55789a  and  a55786a );
 a55791a <=( a55790a  and  a55783a );
 a55794a <=( (not A235)  and  (not A234) );
 a55797a <=( A266  and  A265 );
 a55798a <=( a55797a  and  a55794a );
 a55801a <=( (not A268)  and  (not A267) );
 a55805a <=( (not A302)  and  (not A301) );
 a55806a <=( (not A300)  and  a55805a );
 a55807a <=( a55806a  and  a55801a );
 a55808a <=( a55807a  and  a55798a );
 a55811a <=( (not A169)  and  (not A170) );
 a55814a <=( A199  and  (not A168) );
 a55815a <=( a55814a  and  a55811a );
 a55818a <=( A203  and  (not A200) );
 a55821a <=( A233  and  A232 );
 a55822a <=( a55821a  and  a55818a );
 a55823a <=( a55822a  and  a55815a );
 a55826a <=( (not A235)  and  (not A234) );
 a55829a <=( A266  and  A265 );
 a55830a <=( a55829a  and  a55826a );
 a55833a <=( (not A268)  and  (not A267) );
 a55837a <=( (not A301)  and  (not A299) );
 a55838a <=( (not A298)  and  a55837a );
 a55839a <=( a55838a  and  a55833a );
 a55840a <=( a55839a  and  a55830a );
 a55843a <=( (not A169)  and  (not A170) );
 a55846a <=( A199  and  (not A168) );
 a55847a <=( a55846a  and  a55843a );
 a55850a <=( A203  and  (not A200) );
 a55853a <=( A233  and  A232 );
 a55854a <=( a55853a  and  a55850a );
 a55855a <=( a55854a  and  a55847a );
 a55858a <=( (not A235)  and  (not A234) );
 a55861a <=( (not A266)  and  (not A265) );
 a55862a <=( a55861a  and  a55858a );
 a55865a <=( A298  and  (not A268) );
 a55869a <=( (not A301)  and  (not A300) );
 a55870a <=( A299  and  a55869a );
 a55871a <=( a55870a  and  a55865a );
 a55872a <=( a55871a  and  a55862a );
 a55875a <=( (not A169)  and  (not A170) );
 a55878a <=( A199  and  (not A168) );
 a55879a <=( a55878a  and  a55875a );
 a55882a <=( A203  and  (not A200) );
 a55885a <=( (not A233)  and  (not A232) );
 a55886a <=( a55885a  and  a55882a );
 a55887a <=( a55886a  and  a55879a );
 a55890a <=( A265  and  (not A235) );
 a55893a <=( (not A267)  and  A266 );
 a55894a <=( a55893a  and  a55890a );
 a55897a <=( A298  and  (not A268) );
 a55901a <=( (not A301)  and  (not A300) );
 a55902a <=( A299  and  a55901a );
 a55903a <=( a55902a  and  a55897a );
 a55904a <=( a55903a  and  a55894a );
 a55907a <=( A166  and  A168 );
 a55910a <=( A200  and  A199 );
 a55911a <=( a55910a  and  a55907a );
 a55914a <=( (not A202)  and  (not A201) );
 a55918a <=( (not A234)  and  A233 );
 a55919a <=( A232  and  a55918a );
 a55920a <=( a55919a  and  a55914a );
 a55921a <=( a55920a  and  a55911a );
 a55924a <=( A265  and  (not A235) );
 a55927a <=( (not A267)  and  A266 );
 a55928a <=( a55927a  and  a55924a );
 a55931a <=( A298  and  (not A268) );
 a55935a <=( (not A301)  and  (not A300) );
 a55936a <=( A299  and  a55935a );
 a55937a <=( a55936a  and  a55931a );
 a55938a <=( a55937a  and  a55928a );
 a55941a <=( A167  and  A168 );
 a55944a <=( A200  and  A199 );
 a55945a <=( a55944a  and  a55941a );
 a55948a <=( (not A202)  and  (not A201) );
 a55952a <=( (not A234)  and  A233 );
 a55953a <=( A232  and  a55952a );
 a55954a <=( a55953a  and  a55948a );
 a55955a <=( a55954a  and  a55945a );
 a55958a <=( A265  and  (not A235) );
 a55961a <=( (not A267)  and  A266 );
 a55962a <=( a55961a  and  a55958a );
 a55965a <=( A298  and  (not A268) );
 a55969a <=( (not A301)  and  (not A300) );
 a55970a <=( A299  and  a55969a );
 a55971a <=( a55970a  and  a55965a );
 a55972a <=( a55971a  and  a55962a );
 a55975a <=( A167  and  A170 );
 a55978a <=( (not A201)  and  (not A166) );
 a55979a <=( a55978a  and  a55975a );
 a55982a <=( (not A203)  and  (not A202) );
 a55986a <=( (not A234)  and  A233 );
 a55987a <=( A232  and  a55986a );
 a55988a <=( a55987a  and  a55982a );
 a55989a <=( a55988a  and  a55979a );
 a55992a <=( A265  and  (not A235) );
 a55995a <=( (not A267)  and  A266 );
 a55996a <=( a55995a  and  a55992a );
 a55999a <=( A298  and  (not A268) );
 a56003a <=( (not A301)  and  (not A300) );
 a56004a <=( A299  and  a56003a );
 a56005a <=( a56004a  and  a55999a );
 a56006a <=( a56005a  and  a55996a );
 a56009a <=( A167  and  A170 );
 a56012a <=( A199  and  (not A166) );
 a56013a <=( a56012a  and  a56009a );
 a56016a <=( (not A201)  and  A200 );
 a56020a <=( (not A235)  and  (not A234) );
 a56021a <=( (not A202)  and  a56020a );
 a56022a <=( a56021a  and  a56016a );
 a56023a <=( a56022a  and  a56013a );
 a56026a <=( A265  and  (not A236) );
 a56029a <=( (not A267)  and  A266 );
 a56030a <=( a56029a  and  a56026a );
 a56033a <=( A298  and  (not A268) );
 a56037a <=( (not A301)  and  (not A300) );
 a56038a <=( A299  and  a56037a );
 a56039a <=( a56038a  and  a56033a );
 a56040a <=( a56039a  and  a56030a );
 a56043a <=( A167  and  A170 );
 a56046a <=( A199  and  (not A166) );
 a56047a <=( a56046a  and  a56043a );
 a56050a <=( (not A201)  and  A200 );
 a56054a <=( A233  and  A232 );
 a56055a <=( (not A202)  and  a56054a );
 a56056a <=( a56055a  and  a56050a );
 a56057a <=( a56056a  and  a56047a );
 a56060a <=( (not A235)  and  (not A234) );
 a56063a <=( (not A268)  and  (not A267) );
 a56064a <=( a56063a  and  a56060a );
 a56067a <=( A298  and  (not A269) );
 a56071a <=( (not A301)  and  (not A300) );
 a56072a <=( A299  and  a56071a );
 a56073a <=( a56072a  and  a56067a );
 a56074a <=( a56073a  and  a56064a );
 a56077a <=( A167  and  A170 );
 a56080a <=( A199  and  (not A166) );
 a56081a <=( a56080a  and  a56077a );
 a56084a <=( (not A201)  and  A200 );
 a56088a <=( A233  and  A232 );
 a56089a <=( (not A202)  and  a56088a );
 a56090a <=( a56089a  and  a56084a );
 a56091a <=( a56090a  and  a56081a );
 a56094a <=( (not A235)  and  (not A234) );
 a56097a <=( A266  and  A265 );
 a56098a <=( a56097a  and  a56094a );
 a56101a <=( (not A268)  and  (not A267) );
 a56105a <=( (not A302)  and  (not A301) );
 a56106a <=( (not A300)  and  a56105a );
 a56107a <=( a56106a  and  a56101a );
 a56108a <=( a56107a  and  a56098a );
 a56111a <=( A167  and  A170 );
 a56114a <=( A199  and  (not A166) );
 a56115a <=( a56114a  and  a56111a );
 a56118a <=( (not A201)  and  A200 );
 a56122a <=( A233  and  A232 );
 a56123a <=( (not A202)  and  a56122a );
 a56124a <=( a56123a  and  a56118a );
 a56125a <=( a56124a  and  a56115a );
 a56128a <=( (not A235)  and  (not A234) );
 a56131a <=( A266  and  A265 );
 a56132a <=( a56131a  and  a56128a );
 a56135a <=( (not A268)  and  (not A267) );
 a56139a <=( (not A301)  and  (not A299) );
 a56140a <=( (not A298)  and  a56139a );
 a56141a <=( a56140a  and  a56135a );
 a56142a <=( a56141a  and  a56132a );
 a56145a <=( A167  and  A170 );
 a56148a <=( A199  and  (not A166) );
 a56149a <=( a56148a  and  a56145a );
 a56152a <=( (not A201)  and  A200 );
 a56156a <=( A233  and  A232 );
 a56157a <=( (not A202)  and  a56156a );
 a56158a <=( a56157a  and  a56152a );
 a56159a <=( a56158a  and  a56149a );
 a56162a <=( (not A235)  and  (not A234) );
 a56165a <=( (not A266)  and  (not A265) );
 a56166a <=( a56165a  and  a56162a );
 a56169a <=( A298  and  (not A268) );
 a56173a <=( (not A301)  and  (not A300) );
 a56174a <=( A299  and  a56173a );
 a56175a <=( a56174a  and  a56169a );
 a56176a <=( a56175a  and  a56166a );
 a56179a <=( A167  and  A170 );
 a56182a <=( A199  and  (not A166) );
 a56183a <=( a56182a  and  a56179a );
 a56186a <=( (not A201)  and  A200 );
 a56190a <=( (not A233)  and  (not A232) );
 a56191a <=( (not A202)  and  a56190a );
 a56192a <=( a56191a  and  a56186a );
 a56193a <=( a56192a  and  a56183a );
 a56196a <=( A265  and  (not A235) );
 a56199a <=( (not A267)  and  A266 );
 a56200a <=( a56199a  and  a56196a );
 a56203a <=( A298  and  (not A268) );
 a56207a <=( (not A301)  and  (not A300) );
 a56208a <=( A299  and  a56207a );
 a56209a <=( a56208a  and  a56203a );
 a56210a <=( a56209a  and  a56200a );
 a56213a <=( A167  and  A170 );
 a56216a <=( (not A199)  and  (not A166) );
 a56217a <=( a56216a  and  a56213a );
 a56220a <=( (not A202)  and  (not A200) );
 a56224a <=( (not A234)  and  A233 );
 a56225a <=( A232  and  a56224a );
 a56226a <=( a56225a  and  a56220a );
 a56227a <=( a56226a  and  a56217a );
 a56230a <=( A265  and  (not A235) );
 a56233a <=( (not A267)  and  A266 );
 a56234a <=( a56233a  and  a56230a );
 a56237a <=( A298  and  (not A268) );
 a56241a <=( (not A301)  and  (not A300) );
 a56242a <=( A299  and  a56241a );
 a56243a <=( a56242a  and  a56237a );
 a56244a <=( a56243a  and  a56234a );
 a56247a <=( (not A167)  and  A170 );
 a56250a <=( (not A201)  and  A166 );
 a56251a <=( a56250a  and  a56247a );
 a56254a <=( (not A203)  and  (not A202) );
 a56258a <=( (not A234)  and  A233 );
 a56259a <=( A232  and  a56258a );
 a56260a <=( a56259a  and  a56254a );
 a56261a <=( a56260a  and  a56251a );
 a56264a <=( A265  and  (not A235) );
 a56267a <=( (not A267)  and  A266 );
 a56268a <=( a56267a  and  a56264a );
 a56271a <=( A298  and  (not A268) );
 a56275a <=( (not A301)  and  (not A300) );
 a56276a <=( A299  and  a56275a );
 a56277a <=( a56276a  and  a56271a );
 a56278a <=( a56277a  and  a56268a );
 a56281a <=( (not A167)  and  A170 );
 a56284a <=( A199  and  A166 );
 a56285a <=( a56284a  and  a56281a );
 a56288a <=( (not A201)  and  A200 );
 a56292a <=( (not A235)  and  (not A234) );
 a56293a <=( (not A202)  and  a56292a );
 a56294a <=( a56293a  and  a56288a );
 a56295a <=( a56294a  and  a56285a );
 a56298a <=( A265  and  (not A236) );
 a56301a <=( (not A267)  and  A266 );
 a56302a <=( a56301a  and  a56298a );
 a56305a <=( A298  and  (not A268) );
 a56309a <=( (not A301)  and  (not A300) );
 a56310a <=( A299  and  a56309a );
 a56311a <=( a56310a  and  a56305a );
 a56312a <=( a56311a  and  a56302a );
 a56315a <=( (not A167)  and  A170 );
 a56318a <=( A199  and  A166 );
 a56319a <=( a56318a  and  a56315a );
 a56322a <=( (not A201)  and  A200 );
 a56326a <=( A233  and  A232 );
 a56327a <=( (not A202)  and  a56326a );
 a56328a <=( a56327a  and  a56322a );
 a56329a <=( a56328a  and  a56319a );
 a56332a <=( (not A235)  and  (not A234) );
 a56335a <=( (not A268)  and  (not A267) );
 a56336a <=( a56335a  and  a56332a );
 a56339a <=( A298  and  (not A269) );
 a56343a <=( (not A301)  and  (not A300) );
 a56344a <=( A299  and  a56343a );
 a56345a <=( a56344a  and  a56339a );
 a56346a <=( a56345a  and  a56336a );
 a56349a <=( (not A167)  and  A170 );
 a56352a <=( A199  and  A166 );
 a56353a <=( a56352a  and  a56349a );
 a56356a <=( (not A201)  and  A200 );
 a56360a <=( A233  and  A232 );
 a56361a <=( (not A202)  and  a56360a );
 a56362a <=( a56361a  and  a56356a );
 a56363a <=( a56362a  and  a56353a );
 a56366a <=( (not A235)  and  (not A234) );
 a56369a <=( A266  and  A265 );
 a56370a <=( a56369a  and  a56366a );
 a56373a <=( (not A268)  and  (not A267) );
 a56377a <=( (not A302)  and  (not A301) );
 a56378a <=( (not A300)  and  a56377a );
 a56379a <=( a56378a  and  a56373a );
 a56380a <=( a56379a  and  a56370a );
 a56383a <=( (not A167)  and  A170 );
 a56386a <=( A199  and  A166 );
 a56387a <=( a56386a  and  a56383a );
 a56390a <=( (not A201)  and  A200 );
 a56394a <=( A233  and  A232 );
 a56395a <=( (not A202)  and  a56394a );
 a56396a <=( a56395a  and  a56390a );
 a56397a <=( a56396a  and  a56387a );
 a56400a <=( (not A235)  and  (not A234) );
 a56403a <=( A266  and  A265 );
 a56404a <=( a56403a  and  a56400a );
 a56407a <=( (not A268)  and  (not A267) );
 a56411a <=( (not A301)  and  (not A299) );
 a56412a <=( (not A298)  and  a56411a );
 a56413a <=( a56412a  and  a56407a );
 a56414a <=( a56413a  and  a56404a );
 a56417a <=( (not A167)  and  A170 );
 a56420a <=( A199  and  A166 );
 a56421a <=( a56420a  and  a56417a );
 a56424a <=( (not A201)  and  A200 );
 a56428a <=( A233  and  A232 );
 a56429a <=( (not A202)  and  a56428a );
 a56430a <=( a56429a  and  a56424a );
 a56431a <=( a56430a  and  a56421a );
 a56434a <=( (not A235)  and  (not A234) );
 a56437a <=( (not A266)  and  (not A265) );
 a56438a <=( a56437a  and  a56434a );
 a56441a <=( A298  and  (not A268) );
 a56445a <=( (not A301)  and  (not A300) );
 a56446a <=( A299  and  a56445a );
 a56447a <=( a56446a  and  a56441a );
 a56448a <=( a56447a  and  a56438a );
 a56451a <=( (not A167)  and  A170 );
 a56454a <=( A199  and  A166 );
 a56455a <=( a56454a  and  a56451a );
 a56458a <=( (not A201)  and  A200 );
 a56462a <=( (not A233)  and  (not A232) );
 a56463a <=( (not A202)  and  a56462a );
 a56464a <=( a56463a  and  a56458a );
 a56465a <=( a56464a  and  a56455a );
 a56468a <=( A265  and  (not A235) );
 a56471a <=( (not A267)  and  A266 );
 a56472a <=( a56471a  and  a56468a );
 a56475a <=( A298  and  (not A268) );
 a56479a <=( (not A301)  and  (not A300) );
 a56480a <=( A299  and  a56479a );
 a56481a <=( a56480a  and  a56475a );
 a56482a <=( a56481a  and  a56472a );
 a56485a <=( (not A167)  and  A170 );
 a56488a <=( (not A199)  and  A166 );
 a56489a <=( a56488a  and  a56485a );
 a56492a <=( (not A202)  and  (not A200) );
 a56496a <=( (not A234)  and  A233 );
 a56497a <=( A232  and  a56496a );
 a56498a <=( a56497a  and  a56492a );
 a56499a <=( a56498a  and  a56489a );
 a56502a <=( A265  and  (not A235) );
 a56505a <=( (not A267)  and  A266 );
 a56506a <=( a56505a  and  a56502a );
 a56509a <=( A298  and  (not A268) );
 a56513a <=( (not A301)  and  (not A300) );
 a56514a <=( A299  and  a56513a );
 a56515a <=( a56514a  and  a56509a );
 a56516a <=( a56515a  and  a56506a );
 a56519a <=( (not A167)  and  (not A169) );
 a56522a <=( (not A199)  and  (not A166) );
 a56523a <=( a56522a  and  a56519a );
 a56526a <=( A203  and  A200 );
 a56530a <=( (not A234)  and  A233 );
 a56531a <=( A232  and  a56530a );
 a56532a <=( a56531a  and  a56526a );
 a56533a <=( a56532a  and  a56523a );
 a56536a <=( A265  and  (not A235) );
 a56539a <=( (not A267)  and  A266 );
 a56540a <=( a56539a  and  a56536a );
 a56543a <=( A298  and  (not A268) );
 a56547a <=( (not A301)  and  (not A300) );
 a56548a <=( A299  and  a56547a );
 a56549a <=( a56548a  and  a56543a );
 a56550a <=( a56549a  and  a56540a );
 a56553a <=( (not A167)  and  (not A169) );
 a56556a <=( A199  and  (not A166) );
 a56557a <=( a56556a  and  a56553a );
 a56560a <=( A203  and  (not A200) );
 a56564a <=( (not A234)  and  A233 );
 a56565a <=( A232  and  a56564a );
 a56566a <=( a56565a  and  a56560a );
 a56567a <=( a56566a  and  a56557a );
 a56570a <=( A265  and  (not A235) );
 a56573a <=( (not A267)  and  A266 );
 a56574a <=( a56573a  and  a56570a );
 a56577a <=( A298  and  (not A268) );
 a56581a <=( (not A301)  and  (not A300) );
 a56582a <=( A299  and  a56581a );
 a56583a <=( a56582a  and  a56577a );
 a56584a <=( a56583a  and  a56574a );
 a56587a <=( (not A168)  and  (not A169) );
 a56590a <=( A166  and  A167 );
 a56591a <=( a56590a  and  a56587a );
 a56594a <=( A201  and  A199 );
 a56598a <=( (not A234)  and  A233 );
 a56599a <=( A232  and  a56598a );
 a56600a <=( a56599a  and  a56594a );
 a56601a <=( a56600a  and  a56591a );
 a56604a <=( A265  and  (not A235) );
 a56607a <=( (not A267)  and  A266 );
 a56608a <=( a56607a  and  a56604a );
 a56611a <=( A298  and  (not A268) );
 a56615a <=( (not A301)  and  (not A300) );
 a56616a <=( A299  and  a56615a );
 a56617a <=( a56616a  and  a56611a );
 a56618a <=( a56617a  and  a56608a );
 a56621a <=( (not A168)  and  (not A169) );
 a56624a <=( A166  and  A167 );
 a56625a <=( a56624a  and  a56621a );
 a56628a <=( A201  and  A200 );
 a56632a <=( (not A234)  and  A233 );
 a56633a <=( A232  and  a56632a );
 a56634a <=( a56633a  and  a56628a );
 a56635a <=( a56634a  and  a56625a );
 a56638a <=( A265  and  (not A235) );
 a56641a <=( (not A267)  and  A266 );
 a56642a <=( a56641a  and  a56638a );
 a56645a <=( A298  and  (not A268) );
 a56649a <=( (not A301)  and  (not A300) );
 a56650a <=( A299  and  a56649a );
 a56651a <=( a56650a  and  a56645a );
 a56652a <=( a56651a  and  a56642a );
 a56655a <=( (not A168)  and  (not A169) );
 a56658a <=( A166  and  A167 );
 a56659a <=( a56658a  and  a56655a );
 a56662a <=( A200  and  (not A199) );
 a56666a <=( (not A235)  and  (not A234) );
 a56667a <=( A203  and  a56666a );
 a56668a <=( a56667a  and  a56662a );
 a56669a <=( a56668a  and  a56659a );
 a56672a <=( A265  and  (not A236) );
 a56675a <=( (not A267)  and  A266 );
 a56676a <=( a56675a  and  a56672a );
 a56679a <=( A298  and  (not A268) );
 a56683a <=( (not A301)  and  (not A300) );
 a56684a <=( A299  and  a56683a );
 a56685a <=( a56684a  and  a56679a );
 a56686a <=( a56685a  and  a56676a );
 a56689a <=( (not A168)  and  (not A169) );
 a56692a <=( A166  and  A167 );
 a56693a <=( a56692a  and  a56689a );
 a56696a <=( A200  and  (not A199) );
 a56700a <=( A233  and  A232 );
 a56701a <=( A203  and  a56700a );
 a56702a <=( a56701a  and  a56696a );
 a56703a <=( a56702a  and  a56693a );
 a56706a <=( (not A235)  and  (not A234) );
 a56709a <=( (not A268)  and  (not A267) );
 a56710a <=( a56709a  and  a56706a );
 a56713a <=( A298  and  (not A269) );
 a56717a <=( (not A301)  and  (not A300) );
 a56718a <=( A299  and  a56717a );
 a56719a <=( a56718a  and  a56713a );
 a56720a <=( a56719a  and  a56710a );
 a56723a <=( (not A168)  and  (not A169) );
 a56726a <=( A166  and  A167 );
 a56727a <=( a56726a  and  a56723a );
 a56730a <=( A200  and  (not A199) );
 a56734a <=( A233  and  A232 );
 a56735a <=( A203  and  a56734a );
 a56736a <=( a56735a  and  a56730a );
 a56737a <=( a56736a  and  a56727a );
 a56740a <=( (not A235)  and  (not A234) );
 a56743a <=( A266  and  A265 );
 a56744a <=( a56743a  and  a56740a );
 a56747a <=( (not A268)  and  (not A267) );
 a56751a <=( (not A302)  and  (not A301) );
 a56752a <=( (not A300)  and  a56751a );
 a56753a <=( a56752a  and  a56747a );
 a56754a <=( a56753a  and  a56744a );
 a56757a <=( (not A168)  and  (not A169) );
 a56760a <=( A166  and  A167 );
 a56761a <=( a56760a  and  a56757a );
 a56764a <=( A200  and  (not A199) );
 a56768a <=( A233  and  A232 );
 a56769a <=( A203  and  a56768a );
 a56770a <=( a56769a  and  a56764a );
 a56771a <=( a56770a  and  a56761a );
 a56774a <=( (not A235)  and  (not A234) );
 a56777a <=( A266  and  A265 );
 a56778a <=( a56777a  and  a56774a );
 a56781a <=( (not A268)  and  (not A267) );
 a56785a <=( (not A301)  and  (not A299) );
 a56786a <=( (not A298)  and  a56785a );
 a56787a <=( a56786a  and  a56781a );
 a56788a <=( a56787a  and  a56778a );
 a56791a <=( (not A168)  and  (not A169) );
 a56794a <=( A166  and  A167 );
 a56795a <=( a56794a  and  a56791a );
 a56798a <=( A200  and  (not A199) );
 a56802a <=( A233  and  A232 );
 a56803a <=( A203  and  a56802a );
 a56804a <=( a56803a  and  a56798a );
 a56805a <=( a56804a  and  a56795a );
 a56808a <=( (not A235)  and  (not A234) );
 a56811a <=( (not A266)  and  (not A265) );
 a56812a <=( a56811a  and  a56808a );
 a56815a <=( A298  and  (not A268) );
 a56819a <=( (not A301)  and  (not A300) );
 a56820a <=( A299  and  a56819a );
 a56821a <=( a56820a  and  a56815a );
 a56822a <=( a56821a  and  a56812a );
 a56825a <=( (not A168)  and  (not A169) );
 a56828a <=( A166  and  A167 );
 a56829a <=( a56828a  and  a56825a );
 a56832a <=( A200  and  (not A199) );
 a56836a <=( (not A233)  and  (not A232) );
 a56837a <=( A203  and  a56836a );
 a56838a <=( a56837a  and  a56832a );
 a56839a <=( a56838a  and  a56829a );
 a56842a <=( A265  and  (not A235) );
 a56845a <=( (not A267)  and  A266 );
 a56846a <=( a56845a  and  a56842a );
 a56849a <=( A298  and  (not A268) );
 a56853a <=( (not A301)  and  (not A300) );
 a56854a <=( A299  and  a56853a );
 a56855a <=( a56854a  and  a56849a );
 a56856a <=( a56855a  and  a56846a );
 a56859a <=( (not A168)  and  (not A169) );
 a56862a <=( A166  and  A167 );
 a56863a <=( a56862a  and  a56859a );
 a56866a <=( (not A200)  and  A199 );
 a56870a <=( (not A235)  and  (not A234) );
 a56871a <=( A203  and  a56870a );
 a56872a <=( a56871a  and  a56866a );
 a56873a <=( a56872a  and  a56863a );
 a56876a <=( A265  and  (not A236) );
 a56879a <=( (not A267)  and  A266 );
 a56880a <=( a56879a  and  a56876a );
 a56883a <=( A298  and  (not A268) );
 a56887a <=( (not A301)  and  (not A300) );
 a56888a <=( A299  and  a56887a );
 a56889a <=( a56888a  and  a56883a );
 a56890a <=( a56889a  and  a56880a );
 a56893a <=( (not A168)  and  (not A169) );
 a56896a <=( A166  and  A167 );
 a56897a <=( a56896a  and  a56893a );
 a56900a <=( (not A200)  and  A199 );
 a56904a <=( A233  and  A232 );
 a56905a <=( A203  and  a56904a );
 a56906a <=( a56905a  and  a56900a );
 a56907a <=( a56906a  and  a56897a );
 a56910a <=( (not A235)  and  (not A234) );
 a56913a <=( (not A268)  and  (not A267) );
 a56914a <=( a56913a  and  a56910a );
 a56917a <=( A298  and  (not A269) );
 a56921a <=( (not A301)  and  (not A300) );
 a56922a <=( A299  and  a56921a );
 a56923a <=( a56922a  and  a56917a );
 a56924a <=( a56923a  and  a56914a );
 a56927a <=( (not A168)  and  (not A169) );
 a56930a <=( A166  and  A167 );
 a56931a <=( a56930a  and  a56927a );
 a56934a <=( (not A200)  and  A199 );
 a56938a <=( A233  and  A232 );
 a56939a <=( A203  and  a56938a );
 a56940a <=( a56939a  and  a56934a );
 a56941a <=( a56940a  and  a56931a );
 a56944a <=( (not A235)  and  (not A234) );
 a56947a <=( A266  and  A265 );
 a56948a <=( a56947a  and  a56944a );
 a56951a <=( (not A268)  and  (not A267) );
 a56955a <=( (not A302)  and  (not A301) );
 a56956a <=( (not A300)  and  a56955a );
 a56957a <=( a56956a  and  a56951a );
 a56958a <=( a56957a  and  a56948a );
 a56961a <=( (not A168)  and  (not A169) );
 a56964a <=( A166  and  A167 );
 a56965a <=( a56964a  and  a56961a );
 a56968a <=( (not A200)  and  A199 );
 a56972a <=( A233  and  A232 );
 a56973a <=( A203  and  a56972a );
 a56974a <=( a56973a  and  a56968a );
 a56975a <=( a56974a  and  a56965a );
 a56978a <=( (not A235)  and  (not A234) );
 a56981a <=( A266  and  A265 );
 a56982a <=( a56981a  and  a56978a );
 a56985a <=( (not A268)  and  (not A267) );
 a56989a <=( (not A301)  and  (not A299) );
 a56990a <=( (not A298)  and  a56989a );
 a56991a <=( a56990a  and  a56985a );
 a56992a <=( a56991a  and  a56982a );
 a56995a <=( (not A168)  and  (not A169) );
 a56998a <=( A166  and  A167 );
 a56999a <=( a56998a  and  a56995a );
 a57002a <=( (not A200)  and  A199 );
 a57006a <=( A233  and  A232 );
 a57007a <=( A203  and  a57006a );
 a57008a <=( a57007a  and  a57002a );
 a57009a <=( a57008a  and  a56999a );
 a57012a <=( (not A235)  and  (not A234) );
 a57015a <=( (not A266)  and  (not A265) );
 a57016a <=( a57015a  and  a57012a );
 a57019a <=( A298  and  (not A268) );
 a57023a <=( (not A301)  and  (not A300) );
 a57024a <=( A299  and  a57023a );
 a57025a <=( a57024a  and  a57019a );
 a57026a <=( a57025a  and  a57016a );
 a57029a <=( (not A168)  and  (not A169) );
 a57032a <=( A166  and  A167 );
 a57033a <=( a57032a  and  a57029a );
 a57036a <=( (not A200)  and  A199 );
 a57040a <=( (not A233)  and  (not A232) );
 a57041a <=( A203  and  a57040a );
 a57042a <=( a57041a  and  a57036a );
 a57043a <=( a57042a  and  a57033a );
 a57046a <=( A265  and  (not A235) );
 a57049a <=( (not A267)  and  A266 );
 a57050a <=( a57049a  and  a57046a );
 a57053a <=( A298  and  (not A268) );
 a57057a <=( (not A301)  and  (not A300) );
 a57058a <=( A299  and  a57057a );
 a57059a <=( a57058a  and  a57053a );
 a57060a <=( a57059a  and  a57050a );
 a57063a <=( (not A169)  and  (not A170) );
 a57066a <=( (not A199)  and  (not A168) );
 a57067a <=( a57066a  and  a57063a );
 a57070a <=( A203  and  A200 );
 a57074a <=( (not A234)  and  A233 );
 a57075a <=( A232  and  a57074a );
 a57076a <=( a57075a  and  a57070a );
 a57077a <=( a57076a  and  a57067a );
 a57080a <=( A265  and  (not A235) );
 a57083a <=( (not A267)  and  A266 );
 a57084a <=( a57083a  and  a57080a );
 a57087a <=( A298  and  (not A268) );
 a57091a <=( (not A301)  and  (not A300) );
 a57092a <=( A299  and  a57091a );
 a57093a <=( a57092a  and  a57087a );
 a57094a <=( a57093a  and  a57084a );
 a57097a <=( (not A169)  and  (not A170) );
 a57100a <=( A199  and  (not A168) );
 a57101a <=( a57100a  and  a57097a );
 a57104a <=( A203  and  (not A200) );
 a57108a <=( (not A234)  and  A233 );
 a57109a <=( A232  and  a57108a );
 a57110a <=( a57109a  and  a57104a );
 a57111a <=( a57110a  and  a57101a );
 a57114a <=( A265  and  (not A235) );
 a57117a <=( (not A267)  and  A266 );
 a57118a <=( a57117a  and  a57114a );
 a57121a <=( A298  and  (not A268) );
 a57125a <=( (not A301)  and  (not A300) );
 a57126a <=( A299  and  a57125a );
 a57127a <=( a57126a  and  a57121a );
 a57128a <=( a57127a  and  a57118a );
 a57131a <=( A167  and  A170 );
 a57134a <=( A199  and  (not A166) );
 a57135a <=( a57134a  and  a57131a );
 a57138a <=( (not A201)  and  A200 );
 a57142a <=( A233  and  A232 );
 a57143a <=( (not A202)  and  a57142a );
 a57144a <=( a57143a  and  a57138a );
 a57145a <=( a57144a  and  a57135a );
 a57148a <=( (not A235)  and  (not A234) );
 a57152a <=( (not A267)  and  A266 );
 a57153a <=( A265  and  a57152a );
 a57154a <=( a57153a  and  a57148a );
 a57157a <=( A298  and  (not A268) );
 a57161a <=( (not A301)  and  (not A300) );
 a57162a <=( A299  and  a57161a );
 a57163a <=( a57162a  and  a57157a );
 a57164a <=( a57163a  and  a57154a );
 a57167a <=( (not A167)  and  A170 );
 a57170a <=( A199  and  A166 );
 a57171a <=( a57170a  and  a57167a );
 a57174a <=( (not A201)  and  A200 );
 a57178a <=( A233  and  A232 );
 a57179a <=( (not A202)  and  a57178a );
 a57180a <=( a57179a  and  a57174a );
 a57181a <=( a57180a  and  a57171a );
 a57184a <=( (not A235)  and  (not A234) );
 a57188a <=( (not A267)  and  A266 );
 a57189a <=( A265  and  a57188a );
 a57190a <=( a57189a  and  a57184a );
 a57193a <=( A298  and  (not A268) );
 a57197a <=( (not A301)  and  (not A300) );
 a57198a <=( A299  and  a57197a );
 a57199a <=( a57198a  and  a57193a );
 a57200a <=( a57199a  and  a57190a );
 a57203a <=( (not A168)  and  (not A169) );
 a57206a <=( A166  and  A167 );
 a57207a <=( a57206a  and  a57203a );
 a57210a <=( A200  and  (not A199) );
 a57214a <=( A233  and  A232 );
 a57215a <=( A203  and  a57214a );
 a57216a <=( a57215a  and  a57210a );
 a57217a <=( a57216a  and  a57207a );
 a57220a <=( (not A235)  and  (not A234) );
 a57224a <=( (not A267)  and  A266 );
 a57225a <=( A265  and  a57224a );
 a57226a <=( a57225a  and  a57220a );
 a57229a <=( A298  and  (not A268) );
 a57233a <=( (not A301)  and  (not A300) );
 a57234a <=( A299  and  a57233a );
 a57235a <=( a57234a  and  a57229a );
 a57236a <=( a57235a  and  a57226a );
 a57239a <=( (not A168)  and  (not A169) );
 a57242a <=( A166  and  A167 );
 a57243a <=( a57242a  and  a57239a );
 a57246a <=( (not A200)  and  A199 );
 a57250a <=( A233  and  A232 );
 a57251a <=( A203  and  a57250a );
 a57252a <=( a57251a  and  a57246a );
 a57253a <=( a57252a  and  a57243a );
 a57256a <=( (not A235)  and  (not A234) );
 a57260a <=( (not A267)  and  A266 );
 a57261a <=( A265  and  a57260a );
 a57262a <=( a57261a  and  a57256a );
 a57265a <=( A298  and  (not A268) );
 a57269a <=( (not A301)  and  (not A300) );
 a57270a <=( A299  and  a57269a );
 a57271a <=( a57270a  and  a57265a );
 a57272a <=( a57271a  and  a57262a );


end x25_11x_behav;
